library IEEE;
use IEEE.std_logic_1164.all;

entity somador_tb is
end somador_tb;

architecture arch_somador of somador_tb is

signal clock: std_logic; --:= '0';
signal reset: std_logic; --:= '1'; 
signal wt_in, wt_out: std_logic; 
signal pronto: std_logic; 
signal sela, selb, selc: std_logic; 
signal AB_in, f3_tmp, f3_tmp2, f3, res : std_logic_vector(31 downto 0) := (others => '0');

signal ok, ok_exp, aux: std_logic;
signal auxv1, auxv2 : std_logic_vector(31 downto 0);

type entrada is record
a : std_logic_vector(31 downto 0);
b : std_logic_vector(31 downto 0);
end record;

type test_array is array(positive range <>) of entrada;

	constant test_vector : test_array := (
	(x"00e00000", x"00000000"),
	(x"80800000", x"00600000"),
	(x"00400000", x"00000000"),
	(x"00400000", x"00800000"),
	(x"0980000f", x"00000000"),
	(x"89800000", x"003c0000"),	
	(b"10000000001000010000000000100010", b"00000000000000000000000000000000"),
	(b"10000000001110111001000110100110", b"10000000010111001001000111001000"), -- -3.03062e-39 + -5.47054e-39 = -8.50116e-39
	(b"10000000001010000000100111010100", b"00000000000000000000000000000000"),
	(b"00000000000101101101110010100001", b"10000000000100010010110100110011"), -- -3.67695e-39 + 2.09953e-39 = -1.57742e-39
	(b"00000000001001100011011110111111", b"00000000000000000000000000000000"),
	(b"10000000001000110100000000000110", b"00000000000000101111011110111001"), -- 3.50975e-39 + -3.23721e-39 = 2.72537e-40
	(b"10000000001010101101000000010001", b"00000000000000000000000000000000"),
	(b"00000000001101010100001011010100", b"00000000000010100111001011000011"), -- -3.93173e-39 + 4.89125e-39 = 9.59524e-40
	(b"10000000000101111101010100110010", b"00000000000000000000000000000000"),
	(b"10000000001000011111110111110110", b"10000000001110011101001100101000"), -- -2.1887e-39 + -3.12168e-39 = -5.31037e-39
	(b"00000000001011100111111001100011", b"00000000000000000000000000000000"),
	(b"10000000001111101111101100110101", b"10000000000100000111110011010010"), -- 4.26977e-39 + -5.78392e-39 = -1.51415e-39
	(b"10000000001010010011001100101100", b"00000000000000000000000000000000"),
	(b"10000000001110011010101101110101", b"10000000011000101101111010100001"), -- -3.78361e-39 + -5.29613e-39 = -9.07974e-39
	(b"10000000001101111111110110110001", b"00000000000000000000000000000000"),
	(b"10000000001010011010010000011001", b"10000000011000011010000111001010"), -- -5.14196e-39 + -3.82412e-39 = -8.96608e-39
	(b"10000000000111100100011000101000", b"00000000000000000000000000000000"),
	(b"00000000001101101110011101110111", b"00000000000110001010000101001111"), -- -2.78023e-39 + 5.04215e-39 = 2.26192e-39
	(b"10000000001110000000101000111100", b"00000000000000000000000000000000"),
	(b"00000000000110110110011001001000", b"10000000000111001010001111110100"), -- -5.14646e-39 + 2.51625e-39 = -2.63021e-39
	(b"00000000001101100010000011001011", b"00000000000000000000000000000000"),
	(b"00000000000100001101101000110110", b"00000000010001101111101100000001"), -- 4.97088e-39 + 1.54765e-39 = 6.51853e-39
	(b"00000000001110110010111001001011", b"00000000000000000000000000000000"),
	(b"10000000001011111000000111101000", b"00000000000010111010110001100011"), -- 5.4349e-39 + -4.36287e-39 = 1.07203e-39
	(b"10000000001000011100110100001010", b"00000000000000000000000000000000"),
	(b"00000000001000000011101000111110", b"10000000000000011001001011001100"), -- -3.10413e-39 + 2.95963e-39 = -1.44496e-40
	(b"10000000000111100000010110100000", b"00000000000000000000000000000000"),
	(b"10000000001110001010100001110111", b"10000000010101101010111000010111"), -- -2.75708e-39 + -5.20322e-39 = -7.9603e-39
	(b"10000000000111000110000110101010", b"00000000000000000000000000000000"),
	(b"10000000001011010001111010011100", b"10000000010010011000000001000110"), -- -2.60643e-39 + -4.14358e-39 = -6.75001e-39
	(b"00000000000101100100010100011110", b"00000000000000000000000000000000"),
	(b"10000000000101010101011111011100", b"00000000000000001110110101000010"), -- 2.04518e-39 + -1.96006e-39 = 8.51121e-41
	(b"10000000001011111011010101110011", b"00000000000000000000000000000000"),
	(b"10000000001111001000110001011001", b"10000000011011000100000111001100"), -- -4.38136e-39 + -5.56048e-39 = -9.94184e-39
	(b"00000000001010110010001111101000", b"00000000000000000000000000000000"),
	(b"10000000001111101111100111011011", b"10000000000100111101010111110011"), -- 3.96181e-39 + -5.78343e-39 = -1.82162e-39
	(b"00000000000100100010110111000100", b"00000000000000000000000000000000"),
	(b"10000000001011111111011010011001", b"10000000000111011100100011010101"), -- 1.66946e-39 + -4.40473e-39 = -2.73527e-39
	(b"00000000001011001100101110101110", b"00000000000000000000000000000000"),
	(b"00000000001001110000111011000100", b"00000000010100111101101001110010"), -- 4.11383e-39 + 3.58688e-39 = 7.70071e-39
	(b"00000000001101011110010001010000", b"00000000000000000000000000000000"),
	(b"00000000001101110011100000000000", b"00000000011011010001110001010000"), -- 4.94918e-39 + 5.07104e-39 = 1.00202e-38
	(b"10000000001101101010001001011100", b"00000000000000000000000000000000"),
	(b"00000000000110010001110100000010", b"10000000000111011000010101011010"), -- -5.01736e-39 + 2.30629e-39 = -2.71107e-39
	(b"10000000001001011101101100001110", b"00000000000000000000000000000000"),
	(b"10000000001101011111001101010000", b"10000000010110111100111001011110"), -- -3.4765e-39 + -4.95457e-39 = -8.43106e-39
	(b"00000000001001100101000101001110", b"00000000000000000000000000000000"),
	(b"00000000001111101111001001100001", b"00000000011001010100001110101111"), -- 3.51892e-39 + 5.78075e-39 = 9.29967e-39
	(b"10000000001111010100110011010000", b"00000000000000000000000000000000"),
	(b"10000000001100010100000111110000", b"10000000011011101000111011000000"), -- -5.62952e-39 + -4.52359e-39 = -1.01531e-38
	(b"00000000001011111101111011101101", b"00000000000000000000000000000000"),
	(b"00000000000111001111111111110000", b"00000000010011001101111011011101"), -- 4.39624e-39 + 2.66321e-39 = 7.05945e-39
	(b"10000000000111010100101100000111", b"00000000000000000000000000000000"),
	(b"10000000000110111110011101111110", b"10000000001110010011001010000101"), -- -2.69014e-39 + -2.5626e-39 = -5.25275e-39
	(b"10000000001111100111001010100010", b"00000000000000000000000000000000"),
	(b"10000000000111011011111011011110", b"10000000010111000011000110000000"), -- -5.73492e-39 + -2.7317e-39 = -8.46662e-39
	(b"10000000001000101010111110111111", b"00000000000000000000000000000000"),
	(b"00000000001001011110010001101011", b"00000000000000110011010010101100"), -- -3.18545e-39 + 3.47985e-39 = 2.94402e-40
	(b"00000000001001100110011000000001", b"00000000000000000000000000000000"),
	(b"10000000001000011010001000100111", b"00000000000001001100001111011010"), -- 3.52634e-39 + -3.08874e-39 = 4.376e-40
	(b"00000000000110101001100001111110", b"00000000000000000000000000000000"),
	(b"10000000000101101111110100111101", b"00000000000000111001101101000001"), -- 2.44243e-39 + -2.11123e-39 = 3.31201e-40
	(b"00000000000100000010101011111001", b"00000000000000000000000000000000"),
	(b"10000000000111100100111011011100", b"10000000000011100010001111100011"), -- 1.48478e-39 + -2.78335e-39 = -1.29857e-39
	(b"10000000001110100011000001100111", b"00000000000000000000000000000000"),
	(b"10000000001000011000111111001101", b"10000000010110111100000000110100"), -- -5.34382e-39 + -3.08216e-39 = -8.42598e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011111110010000000110011", b"11111111100000000000000000000000"), -- -inf + 1.16747e-38 = -inf
	(b"00111010001010010001110111010101", b"00000000000000000000000000000000"),
	(b"10000000000011101110011001110111", b"00111010001010010001110111010101"), -- 0.000645128 + -1.36837e-39 = 0.000645128
	(b"11001101110010111011000000001101", b"00000000000000000000000000000000"),
	(b"00000000011010000111110110100001", b"11001101110010111011000000001101"), -- -4.27164e+08 + 9.59596e-39 = -4.27164e+08
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110110011100101001000", b"10000000011110110011100101001000"), -- 0 + -1.13163e-38 = -1.13163e-38
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000111111100001001110", b"10000000000000111111100001001110"), -- 0 + -3.64581e-40 = -3.64581e-40
	(b"00000000000000000000000010000110", b"00000000000000000000000000000000"),
	(b"10000000001101110100111111110101", b"10000000001101110100111101101111"), -- 1.87774e-43 + -5.07964e-39 = -5.07945e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001111111100101101111", b"01111111100000000000000000000000"), -- inf + -3.67106e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110000111011010000011", b"01111111100000000000000000000000"), -- inf + 8.12404e-39 = inf
	(b"11011001110111101010001010001100", b"00000000000000000000000000000000"),
	(b"10000000011001101110110010111010", b"11011001110111101010001010001100"), -- -7.83327e+15 + -9.45214e-39 = -7.83327e+15
	(b"00111000100011110010101101010111", b"00000000000000000000000000000000"),
	(b"00000000011011100011100111110111", b"00111000100011110010101101010111"), -- 6.82684e-05 + 1.01227e-38 = 6.82684e-05
	(b"11011000001101011001110101001111", b"00000000000000000000000000000000"),
	(b"00000000000010111000010110011101", b"11011000001101011001110101001111"), -- -7.98749e+14 + 1.05812e-39 = -7.98749e+14
	(b"00001000011110111111001110010101", b"00000000000000000000000000000000"),
	(b"00000000000011010111001110001001", b"00001000011110111111001110110000"), -- 7.58189e-34 + 1.23531e-39 = 7.5819e-34
	(b"01010100111100100000101001011010", b"00000000000000000000000000000000"),
	(b"00000000001110000111011001001000", b"01010100111100100000101001011010"), -- 8.31645e+12 + 5.18522e-39 = 8.31645e+12
	(b"10111000101111001101011100100111", b"00000000000000000000000000000000"),
	(b"10000000001001100111101011101110", b"10111000101111001101011100100111"), -- -9.00461e-05 + -3.53385e-39 = -9.00461e-05
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001101000110110100100", b"00000000011001101000110110100100"), -- -0 + 9.41803e-39 = 9.41803e-39
	(b"11010110011011010001100011101001", b"00000000000000000000000000000000"),
	(b"00000000011100101001111100101000", b"11010110011011010001100011101001"), -- -6.51728e+13 + 1.05263e-38 = -6.51728e+13
	(b"10010100010111110011010010100010", b"00000000000000000000000000000000"),
	(b"00000000000011000110001101001111", b"10010100010111110011010010100010"), -- -1.1269e-26 + 1.13765e-39 = -1.1269e-26
	(b"11010100011111111111001100010010", b"00000000000000000000000000000000"),
	(b"00000000001101101110101100001100", b"11010100011111111111001100010010"), -- -4.39718e+12 + 5.04344e-39 = -4.39718e+12
	(b"10111111111000001011110000101110", b"00000000000000000000000000000000"),
	(b"00000000000101111000111110001101", b"10111111111000001011110000101110"), -- -1.75574 + 2.16371e-39 = -1.75574
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011010011111111001001", b"11111111100000000000000000000000"), -- -inf + 4.15548e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010100110100111110001000", b"11111111100000000000000000000000"), -- -inf + 7.65088e-39 = -inf
	(b"10110111110110101101100110010100", b"00000000000000000000000000000000"),
	(b"10000000000011001011111110010011", b"10110111110110101101100110010100"), -- -2.60889e-05 + -1.17075e-39 = -2.60889e-05
	(b"01011000100010011110111110101111", b"00000000000000000000000000000000"),
	(b"10000000010100010101000001011100", b"01011000100010011110111110101111"), -- 1.2133e+15 + -7.4675e-39 = 1.2133e+15
	(b"01101110100010010000011010101111", b"00000000000000000000000000000000"),
	(b"10000000010110001011001110000000", b"01101110100010010000011010101111"), -- 2.12038e+28 + -8.14592e-39 = 2.12038e+28
	(b"10101110000011110101000011111100", b"00000000000000000000000000000000"),
	(b"00000000000100011010010000110101", b"10101110000011110101000011111100"), -- -3.25864e-11 + 1.62011e-39 = -3.25864e-11
	(b"00100001001100101011010110101010", b"00000000000000000000000000000000"),
	(b"10000000010110011011011110011110", b"00100001001100101011010110101010"), -- 6.05492e-19 + -8.23923e-39 = 6.05492e-19
	(b"00011110111100001100101111110010", b"00000000000000000000000000000000"),
	(b"10000000010011000010111101000011", b"00011110111100001100101111110010"), -- 2.54953e-20 + -6.99645e-39 = 2.54953e-20
	(b"10000000000000000000000001100010", b"00000000000000000000000000000000"),
	(b"00000000000001101000111100011010", b"00000000000001101000111010111000"), -- -1.37327e-43 + 6.02348e-40 = 6.02211e-40
	(b"11000100011010010010111010001011", b"00000000000000000000000000000000"),
	(b"00000000001110010111100101001001", b"11000100011010010010111010001011"), -- -932.727 + 5.27813e-39 = -932.727
	(b"10000001110011111010110010101110", b"00000000000000000000000000000000"),
	(b"00000000001000011100011110111101", b"10000001110001110011101010111111"), -- -7.62876e-38 + 3.10222e-39 = -7.31854e-38
	(b"00110001101111110100101011001001", b"00000000000000000000000000000000"),
	(b"00000000001100111011011000110110", b"00110001101111110100101011001001"), -- 5.56733e-09 + 4.74898e-39 = 5.56733e-09
	(b"01011111111111101110000101001011", b"00000000000000000000000000000000"),
	(b"00000000010010101110010010100111", b"01011111111111101110000101001011"), -- 3.67321e+19 + 6.87785e-39 = 3.67321e+19
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011111011111100011101", b"01111111100000000000000000000000"), -- inf + 1.44609e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001101100000010010001", b"00000000000001101100000010010001"), -- 0 + 6.20093e-40 = 6.20093e-40
	(b"10001011000010001000010111111110", b"00000000000000000000000000000000"),
	(b"00000000010101000101010000100110", b"10001011000010001000010111111011"), -- -2.62935e-32 + 7.74437e-39 = -2.62934e-32
	(b"11000010100001100011100000010000", b"00000000000000000000000000000000"),
	(b"00000000011110110001010011001111", b"11000010100001100011100000010000"), -- -67.1095 + 1.13032e-38 = -67.1095
	(b"11101001011110101010011101100001", b"00000000000000000000000000000000"),
	(b"10000000001000010010011100110111", b"11101001011110101010011101100001"), -- -1.89389e+25 + -3.04464e-39 = -1.89389e+25
	(b"01000110000101100011001100111100", b"00000000000000000000000000000000"),
	(b"00000000011100100011001000001000", b"01000110000101100011001100111100"), -- 9612.81 + 1.04872e-38 = 9612.81
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001111010010110001001110", b"01111111100000000000000000000000"), -- inf + -5.61786e-39 = inf
	(b"11000101010000110001010111110110", b"00000000000000000000000000000000"),
	(b"00000000011110100000100010011000", b"11000101010000110001010111110110"), -- -3121.37 + 1.1207e-38 = -3121.37
	(b"00001110111000000101100000101101", b"00000000000000000000000000000000"),
	(b"10000000000011111011110011100000", b"00001110111000000101100000101101"), -- 5.53052e-30 + -1.44529e-39 = 5.53052e-30
	(b"10111000110101101001011010001111", b"00000000000000000000000000000000"),
	(b"00000000000001011110101000000000", b"10111000110101101001011010001111"), -- -0.000102324 + 5.43121e-40 = -0.000102324
	(b"00111100001011110001110100001001", b"00000000000000000000000000000000"),
	(b"10000000010001101100101010110101", b"00111100001011110001110100001001"), -- 0.0106881 + -6.5012e-39 = 0.0106881
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000101001011010000100111", b"01111111100000000000000000000000"), -- inf + -1.90134e-39 = inf
	(b"00110111010010011001111111010001", b"00000000000000000000000000000000"),
	(b"10000000000101010101010011110110", b"00110111010010011001111111010001"), -- 1.20177e-05 + -1.95902e-39 = 1.20177e-05
	(b"01111100110111010000001001011110", b"00000000000000000000000000000000"),
	(b"10000000001000000110111011101000", b"01111100110111010000001001011110"), -- 9.18036e+36 + -2.97852e-39 = 9.18036e+36
	(b"11101111100000011000000010111111", b"00000000000000000000000000000000"),
	(b"00000000010010000001100101111000", b"11101111100000011000000010111111"), -- -8.01584e+28 + 6.62129e-39 = -8.01584e+28
	(b"11000011011000101001011111001101", b"00000000000000000000000000000000"),
	(b"00000000001100000100000001001001", b"11000011011000101001011111001101"), -- -226.593 + 4.43116e-39 = -226.593
	(b"00110100010010011011000110100011", b"00000000000000000000000000000000"),
	(b"10000000011011100100101111101011", b"00110100010010011011000110100011"), -- 1.87842e-07 + -1.01291e-38 = 1.87842e-07
	(b"10100110001000001100111101001100", b"00000000000000000000000000000000"),
	(b"10000000000110011010111011001101", b"10100110001000001100111101001100"), -- -5.57921e-16 + -2.35859e-39 = -5.57921e-16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000101001100001001010110", b"10000000000101001100001001010110"), -- 0 + -1.90642e-39 = -1.90642e-39
	(b"01000111110111000100110110111010", b"00000000000000000000000000000000"),
	(b"00000000010101101110101111110111", b"01000111110111000100110110111010"), -- 112795 + 7.9825e-39 = 112795
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000110101111111001010", b"00000000001000110101111111001010"), -- -0 + 3.24861e-39 = 3.24861e-39
	(b"10000000111010111110110001101111", b"00000000000000000000000000000000"),
	(b"10000000001110110111001110010000", b"10000001000100111011000000000000"), -- -2.16662e-38 + -5.45975e-39 = -2.71259e-38
	(b"01000000110010010101110101101111", b"00000000000000000000000000000000"),
	(b"00000000000110001011010000000110", b"01000000110010010101110101101111"), -- 6.29266 + 2.26863e-39 = 6.29266
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010100110011110010101110", b"00000000010100110011110010101110"), -- -0 + 7.64411e-39 = 7.64411e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000111011001110011101", b"01111111100000000000000000000000"), -- inf + -3.3994e-40 = inf
	(b"10100110110101011010100111110100", b"00000000000000000000000000000000"),
	(b"10000000011010110010100110011000", b"10100110110101011010100111110100"), -- -1.48259e-15 + -9.84132e-39 = -1.48259e-15
	(b"00100101010010000000001000000110", b"00000000000000000000000000000000"),
	(b"00000000000010111100100100111011", b"00100101010010000000001000000110"), -- 1.73479e-16 + 1.08238e-39 = 1.73479e-16
	(b"01010000100110111010100100011001", b"00000000000000000000000000000000"),
	(b"00000000000000011110000110100001", b"01010000100110111010100100011001"), -- 2.08924e+10 + 1.72776e-40 = 2.08924e+10
	(b"01110111010010010001001110001000", b"00000000000000000000000000000000"),
	(b"00000000000111100111010111011001", b"01110111010010010001001110001000"), -- 4.07831e+33 + 2.79734e-39 = 4.07831e+33
	(b"01001110101011000100101001101000", b"00000000000000000000000000000000"),
	(b"10000000011100011100110110101011", b"01001110101011000100101001101000"), -- 1.44528e+09 + -1.04512e-38 = 1.44528e+09
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110001010101101110111", b"00000000000110001010101101110111"), -- 0 + 2.26556e-39 = 2.26556e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010100010001101011000101", b"10000000010100010001101011000101"), -- 0 + -7.44828e-39 = -7.44828e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001101100011000110010", b"00000000010001101100011000110010"), -- 0 + 6.49958e-39 = 6.49958e-39
	(b"00111001100011110111001011101101", b"00000000000000000000000000000000"),
	(b"00000000010010011001001110110001", b"00111001100011110111001011101101"), -- 0.000273607 + 6.75697e-39 = 0.000273607
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001100110111110010101010", b"00000000001100110111110010101010"), -- -0 + 4.72833e-39 = 4.72833e-39
	(b"10101011011011110000000001110010", b"00000000000000000000000000000000"),
	(b"10000000011111100110100001100001", b"10101011011011110000000001110010"), -- -8.49105e-13 + -1.16087e-38 = -8.49105e-13
	(b"10000000000000000000000001101100", b"00000000000000000000000000000000"),
	(b"00000000010101111111101000100100", b"00000000010101111111100110111000"), -- -1.5134e-43 + 8.07942e-39 = 8.07927e-39
	(b"00100101001000111010110111000110", b"00000000000000000000000000000000"),
	(b"10000000001001001001001111100010", b"00100101001000111010110111000110"), -- 1.41969e-16 + -3.35913e-39 = 1.41969e-16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110000101101100010011", b"01111111100000000000000000000000"), -- inf + 8.11419e-39 = inf
	(b"01010001101001110100111000010010", b"00000000000000000000000000000000"),
	(b"00000000000101000101111101110110", b"01010001101001110100111000010010"), -- 8.98212e+10 + 1.87095e-39 = 8.98212e+10
	(b"00001101010001011110101000100110", b"00000000000000000000000000000000"),
	(b"00000000000001001110011011101101", b"00001101010001011110101000100110"), -- 6.09872e-31 + 4.50183e-40 = 6.09872e-31
	(b"01011000110000110110010110001100", b"00000000000000000000000000000000"),
	(b"10000000000101110000000011000111", b"01011000110000110110010110001100"), -- 1.71873e+15 + -2.1125e-39 = 1.71873e+15
	(b"01101000111000111010010000111100", b"00000000000000000000000000000000"),
	(b"00000000000011100001101010111000", b"01101000111000111010010000111100"), -- 8.60005e+24 + 1.29528e-39 = 8.60005e+24
	(b"00100111001101010110110100111000", b"00000000000000000000000000000000"),
	(b"00000000010100010101010010110000", b"00100111001101010110110100111000"), -- 2.5178e-15 + 7.46906e-39 = 2.5178e-15
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010000111100101110110100", b"11111111100000000000000000000000"), -- -inf + -6.22605e-39 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010010010000100000110", b"10000000001010010010000100000110"), -- 0 + -3.7771e-39 = -3.7771e-39
	(b"10010000010001110000111011001010", b"00000000000000000000000000000000"),
	(b"00000000011100110110000100111000", b"10010000010001110000111011001010"), -- -3.92572e-29 + 1.0596e-38 = -3.92572e-29
	(b"10111100011100111101010110111101", b"00000000000000000000000000000000"),
	(b"10000000001011101001101010101000", b"10111100011100111101010110111101"), -- -0.0148825 + -4.27991e-39 = -0.0148825
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011110001011100100011", b"10000000000011110001011100100011"), -- 0 + -1.38583e-39 = -1.38583e-39
	(b"11001000001001011001000101100101", b"00000000000000000000000000000000"),
	(b"00000000000010111010101110000001", b"11001000001001011001000101100101"), -- -169542 + 1.07171e-39 = -169542
	(b"10011011001100100100010011001101", b"00000000000000000000000000000000"),
	(b"00000000010110001000000011101101", b"10011011001100100100010011001101"), -- -1.4746e-22 + 8.12777e-39 = -1.4746e-22
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110100100010001110101", b"10000000010110100100010001110101"), -- 0 + -8.28975e-39 = -8.28975e-39
	(b"10011000001010100010101011101110", b"00000000000000000000000000000000"),
	(b"10000000011000111101011100010101", b"10011000001010100010101011101110"), -- -2.19937e-24 + -9.16887e-39 = -2.19937e-24
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011100011011100100010", b"01111111100000000000000000000000"), -- inf + 4.24421e-39 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101101111110110111100", b"10000000011101101111110110111100"), -- -0 + -1.09276e-38 = -1.09276e-38
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100110001100000010100", b"10000000000100110001100000010100"), -- -0 + -1.75351e-39 = -1.75351e-39
	(b"11011110100101001100110111110111", b"00000000000000000000000000000000"),
	(b"00000000010111101100111000010100", b"11011110100101001100110111110111"), -- -5.36125e+18 + 8.70646e-39 = -5.36125e+18
	(b"01001110011010111110101001110111", b"00000000000000000000000000000000"),
	(b"00000000010010101010110101001011", b"01001110011010111110101001110111"), -- 9.89503e+08 + 6.85799e-39 = 9.89503e+08
	(b"00110110010110101010000001101001", b"00000000000000000000000000000000"),
	(b"10000000010000001000011000100111", b"00110110010110101010000001101001"), -- 3.25779e-06 + -5.9256e-39 = 3.25779e-06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011111000111000100101", b"00000000000011111000111000100101"), -- 0 + 1.42852e-39 = 1.42852e-39
	(b"00100100011001000111010010001000", b"00000000000000000000000000000000"),
	(b"00000000001110000011100100011100", b"00100100011001000111010010001000"), -- 4.95383e-17 + 5.16327e-39 = 4.95383e-17
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101110111111100010100", b"01111111100000000000000000000000"), -- inf + 1.0974e-38 = inf
	(b"10111010111010000100010100000110", b"00000000000000000000000000000000"),
	(b"00000000010101101000010111100010", b"10111010111010000100010100000110"), -- -0.00177208 + 7.94588e-39 = -0.00177208
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111100101101001101110", b"01111111100000000000000000000000"), -- inf + 5.72624e-39 = inf
	(b"11001010111110010110110001111001", b"00000000000000000000000000000000"),
	(b"00000000000000101000000110010000", b"11001010111110010110110001111001"), -- -8.17312e+06 + 2.30149e-40 = -8.17312e+06
	(b"10110110100100101101100110110110", b"00000000000000000000000000000000"),
	(b"00000000010011011111010101010101", b"10110110100100101101100110110110"), -- -4.37648e-06 + 7.15934e-39 = -4.37648e-06
	(b"11110010110000111001111101001110", b"00000000000000000000000000000000"),
	(b"10000000000100001000111011011111", b"11110010110000111001111101001110"), -- -7.7494e+30 + -1.52062e-39 = -7.7494e+30
	(b"00011010011001010000101101101101", b"00000000000000000000000000000000"),
	(b"00000000001111100010101011010101", b"00011010011001010000101101101101"), -- 4.73653e-23 + 5.70917e-39 = 4.73653e-23
	(b"01100111100011000101011100000110", b"00000000000000000000000000000000"),
	(b"10000000000111001101011101101111", b"01100111100011000101011100000110"), -- 1.32547e+24 + -2.64868e-39 = 1.32547e+24
	(b"01011011101101111000110110011000", b"00000000000000000000000000000000"),
	(b"10000000001010110110101001011011", b"01011011101101111000110110011000"), -- 1.03331e+17 + -3.98708e-39 = 1.03331e+17
	(b"11000011111001101101011001100100", b"00000000000000000000000000000000"),
	(b"00000000001110010010000000000011", b"11000011111001101101011001100100"), -- -461.675 + 5.24611e-39 = -461.675
	(b"00011011001100001100000000100111", b"00000000000000000000000000000000"),
	(b"00000000000101010101100010000110", b"00011011001100001100000000100111"), -- 1.46205e-22 + 1.9603e-39 = 1.46205e-22
	(b"01000101011111011111010001111011", b"00000000000000000000000000000000"),
	(b"10000000001111101110110101110101", b"01000101011111011111010001111011"), -- 4063.28 + -5.77898e-39 = 4063.28
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001001100111001000000001", b"11111111100000000000000000000000"), -- -inf + 3.53065e-39 = -inf
	(b"11001001111111100101101010000101", b"00000000000000000000000000000000"),
	(b"00000000011011111001101100001111", b"11001001111111100101101010000101"), -- -2.08366e+06 + 1.02494e-38 = -2.08366e+06
	(b"01000010000011100101001011001001", b"00000000000000000000000000000000"),
	(b"00000000000001010001111011010110", b"01000010000011100101001011001001"), -- 35.5808 + 4.70239e-40 = 35.5808
	(b"01001011110100101000100010100110", b"00000000000000000000000000000000"),
	(b"10000000001100001101011000011110", b"01001011110100101000100010100110"), -- 2.75951e+07 + -4.48491e-39 = 2.75951e+07
	(b"10011000000000110011110001011111", b"00000000000000000000000000000000"),
	(b"10000000000101111110010010101000", b"10011000000000110011110001011111"), -- -1.69618e-24 + -2.19424e-39 = -1.69618e-24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001101011111010001011110", b"00000000001101011111010001011110"), -- -0 + 4.95494e-39 = 4.95494e-39
	(b"10101100101111111010101000011011", b"00000000000000000000000000000000"),
	(b"00000000010001111111001111000111", b"10101100101111111010101000011011"), -- -5.44743e-12 + 6.60777e-39 = -5.44743e-12
	(b"01100110101011011001000100101111", b"00000000000000000000000000000000"),
	(b"00000000001100000000010001000001", b"01100110101011011001000100101111"), -- 4.09824e+23 + 4.40963e-39 = 4.09824e+23
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011000111111101000010", b"00000000000011000111111101000010"), -- -0 + 1.14768e-39 = 1.14768e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101111010100011010110", b"10000000011101111010100011010110"), -- 0 + -1.0989e-38 = -1.0989e-38
	(b"01101001010010110000011101101110", b"00000000000000000000000000000000"),
	(b"00000000001010010101101100011000", b"01101001010010110000011101101110"), -- 1.53404e+25 + 3.79793e-39 = 1.53404e+25
	(b"00000000000000000010010101000011", b"00000000000000000000000000000000"),
	(b"00000000000100011001100010101101", b"00000000000100011011110111110000"), -- 1.3367e-41 + 1.61597e-39 = 1.62934e-39
	(b"01111001000111011001000010001011", b"00000000000000000000000000000000"),
	(b"00000000010001000000000000111010", b"01111001000111011001000010001011"), -- 5.11326e+34 + 6.2449e-39 = 5.11326e+34
	(b"00100101100000001110110001101000", b"00000000000000000000000000000000"),
	(b"10000000001100100000111011111001", b"00100101100000001110110001101000"), -- 2.23647e-16 + -4.59715e-39 = 2.23647e-16
	(b"00111110000011110101011101100000", b"00000000000000000000000000000000"),
	(b"10000000010110101010011011110100", b"00111110000011110101011101100000"), -- 0.139982 + -8.32509e-39 = 0.139982
	(b"01101101001100111110011100001110", b"00000000000000000000000000000000"),
	(b"00000000011101110010001100010110", b"01101101001100111110011100001110"), -- 3.47982e+27 + 1.0941e-38 = 3.47982e+27
	(b"00011110010100101100110100101100", b"00000000000000000000000000000000"),
	(b"10000000000100101111111011001111", b"00011110010100101100110100101100"), -- 1.11597e-20 + -1.74445e-39 = 1.11597e-20
	(b"01011101011011011010101011100111", b"00000000000000000000000000000000"),
	(b"10000000000011110110000001010111", b"01011101011011011010101011100111"), -- 1.07036e+18 + -1.41209e-39 = 1.07036e+18
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110001111000111010111", b"00000000000110001111000111010111"), -- 0 + 2.29081e-39 = 2.29081e-39
	(b"11010100011000111100000010101010", b"00000000000000000000000000000000"),
	(b"00000000001100111111110111110000", b"11010100011000111100000010101010"), -- -3.91276e+12 + 4.77471e-39 = -3.91276e+12
	(b"11100101011000110110001100001101", b"00000000000000000000000000000000"),
	(b"10000000001100101110000111001101", b"11100101011000110110001100001101"), -- -6.71128e+22 + -4.67278e-39 = -6.71128e+22
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000001111110000111101111", b"10000000000001111110000111101111"), -- 0 + -7.23898e-40 = -7.23898e-40
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010011001001101101100", b"00000000001010011001001101101100"), -- 0 + 3.81814e-39 = 3.81814e-39
	(b"10001101101111000100100111100111", b"00000000000000000000000000000000"),
	(b"10000000000001100010101000111011", b"10001101101111000100100111100111"), -- -1.16042e-30 + -5.66162e-40 = -1.16042e-30
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001000101010100100000", b"11111111100000000000000000000000"), -- -inf + -3.33661e-39 = -inf
	(b"10001000011011011011111011001001", b"00000000000000000000000000000000"),
	(b"00000000011110100011010010100111", b"10001000011011011011110111010101"), -- -7.15439e-34 + 1.12228e-38 = -7.15427e-34
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001010100011000011111", b"11111111100000000000000000000000"), -- -inf + -9.30054e-39 = -inf
	(b"00101101100001010010111111100011", b"00000000000000000000000000000000"),
	(b"00000000001101110011010000100000", b"00101101100001010010111111100011"), -- 1.51416e-11 + 5.06965e-39 = 1.51416e-11
	(b"00011000010110110011010101011100", b"00000000000000000000000000000000"),
	(b"00000000011100100101101101110111", b"00011000010110110011010101011100"), -- 2.8332e-24 + 1.05021e-38 = 2.8332e-24
	(b"00000000000000000000000000001010", b"00000000000000000000000000000000"),
	(b"10000000010001001100100111110101", b"10000000010001001100100111101011"), -- 1.4013e-44 + -6.31726e-39 = -6.31725e-39
	(b"00001011001001000010110111101011", b"00000000000000000000000000000000"),
	(b"00000000011000110011001101100100", b"00001011001001000010110111101110"), -- 3.16198e-32 + 9.11015e-39 = 3.16198e-32
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011111110101101110111", b"00000000000011111110101101110111"), -- -0 + 1.462e-39 = 1.462e-39
	(b"01001110110111100100110000000110", b"00000000000000000000000000000000"),
	(b"10000000011011111111001111101100", b"01001110110111100100110000000110"), -- 1.86476e+09 + -1.02812e-38 = 1.86476e+09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001010011110111100100", b"01111111100000000000000000000000"), -- inf + 9.29759e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000110001110011110011", b"11111111100000000000000000000000"), -- -inf + -9.1021e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011010000101100101000", b"11111111100000000000000000000000"), -- -inf + -1.19786e-39 = -inf
	(b"10010111100111111110001010101011", b"00000000000000000000000000000000"),
	(b"00000000011100101000011000101001", b"10010111100111111110001010101011"), -- -1.03324e-24 + 1.05174e-38 = -1.03324e-24
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010001101101000111010001", b"01111111100000000000000000000000"), -- inf + -6.50375e-39 = inf
	(b"11011000001110000001000010010000", b"00000000000000000000000000000000"),
	(b"10000000010000110100111100101000", b"11011000001110000001000010010000"), -- -8.09525e+14 + -6.18137e-39 = -8.09525e+14
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111001110101001110111", b"00000000000111001110101001110111"), -- 0 + 2.6555e-39 = 2.6555e-39
	(b"11001001000000001001101100010010", b"00000000000000000000000000000000"),
	(b"00000000011110101111110100000000", b"11001001000000001001101100010010"), -- -526769 + 1.12947e-38 = -526769
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000001100011010000100", b"11111111100000000000000000000000"), -- -inf + 7.1214e-41 = -inf
	(b"10011101000011011000110010110000", b"00000000000000000000000000000000"),
	(b"10000000000110100000011011110101", b"10011101000011011000110010110000"), -- -1.87339e-21 + -2.39022e-39 = -1.87339e-21
	(b"00010111110110111011100010011011", b"00000000000000000000000000000000"),
	(b"00000000000101000000011101111100", b"00010111110110111011100010011011"), -- 1.41991e-24 + 1.83939e-39 = 1.41991e-24
	(b"01010101010000100010010000111000", b"00000000000000000000000000000000"),
	(b"10000000010000001001011011100111", b"01010101010000100010010000111000"), -- 1.33413e+13 + -5.93161e-39 = 1.33413e+13
	(b"01100000100010001100001010110100", b"00000000000000000000000000000000"),
	(b"10000000011011111010100101100100", b"01100000100010001100001010110100"), -- 7.88371e+19 + -1.02545e-38 = 7.88371e+19
	(b"00000000000011001011100101011100", b"00000000000000000000000000000000"),
	(b"00000000010000010001101001111000", b"00000000010011011101001111010100"), -- 1.16852e-39 + 5.9788e-39 = 7.14732e-39
	(b"00110100101010000010101111000111", b"00000000000000000000000000000000"),
	(b"10000000011111010101110110101111", b"00110100101010000010101111000111"), -- 3.13243e-07 + -1.1513e-38 = 3.13243e-07
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110101011100110011111", b"01111111100000000000000000000000"), -- inf + 5.39305e-39 = inf
	(b"11010000100110101000010000110000", b"00000000000000000000000000000000"),
	(b"00000000011101101010011110010100", b"11010000100110101000010000110000"), -- -2.07388e+10 + 1.08967e-38 = -2.07388e+10
	(b"10000000000000000000000110101111", b"00000000000000000000000000000000"),
	(b"00000000001000000001010000100010", b"00000000001000000001001001110011"), -- -6.0396e-43 + 2.94596e-39 = 2.94535e-39
	(b"01000001110001111110011011001101", b"00000000000000000000000000000000"),
	(b"10000000010000100110101111100000", b"01000001110001111110011011001101"), -- 24.9877 + -6.09984e-39 = 24.9877
	(b"11010001010011100100111010101010", b"00000000000000000000000000000000"),
	(b"10000000000011101111101011001100", b"11010001010011100100111010101010"), -- -5.53802e+10 + -1.37567e-39 = -5.53802e+10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010011001010010000010", b"11111111100000000000000000000000"), -- -inf + 8.79794e-40 = -inf
	(b"10000000000000000000000001111010", b"00000000000000000000000000000000"),
	(b"10000000000110101010001001000101", b"10000000000110101010001010111111"), -- -1.70958e-43 + -2.44593e-39 = -2.44611e-39
	(b"00110101010000000000111101000010", b"00000000000000000000000000000000"),
	(b"10000000011111110010000011001011", b"00110101010000000000111101000010"), -- 7.15478e-07 + -1.16749e-38 = 7.15478e-07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010010101110011011010", b"00000000000010010101110011011010"), -- -0 + 8.59828e-40 = 8.59828e-40
	(b"11111010010011000001111101100110", b"00000000000000000000000000000000"),
	(b"00000000000001000000110111110000", b"11111010010011000001111101100110"), -- -2.64966e+35 + 3.72342e-40 = -2.64966e+35
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100100010000001110011", b"01111111100000000000000000000000"), -- inf + 1.66468e-39 = inf
	(b"11000000110100100101101100011000", b"00000000000000000000000000000000"),
	(b"00000000011001000000101111100001", b"11000000110100100101101100011000"), -- -6.57362 + 9.18781e-39 = -6.57362
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010000001110101100000100", b"10000000010000001110101100000100"), -- 0 + -5.96178e-39 = -5.96178e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100101001010100010101", b"11111111100000000000000000000000"), -- -inf + 1.70652e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001111011010110111111111", b"11111111100000000000000000000000"), -- -inf + -5.66438e-39 = -inf
	(b"11010101000011011001001010100100", b"00000000000000000000000000000000"),
	(b"10000000011110110111000110110100", b"11010101000011011001001010100100"), -- -9.72881e+12 + -1.13366e-38 = -9.72881e+12
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010011100111001010110", b"01111111100000000000000000000000"), -- inf + 3.83927e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001011101111011110111", b"11111111100000000000000000000000"), -- -inf + 9.35537e-39 = -inf
	(b"01110111000111011011101111100001", b"00000000000000000000000000000000"),
	(b"00000000000011011100011010001110", b"01110111000111011011101111100001"), -- 3.19922e+33 + 1.26509e-39 = 3.19922e+33
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011010100001000001001011", b"01111111100000000000000000000000"), -- inf + 9.74041e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010010011011001111100", b"01111111100000000000000000000000"), -- inf + -3.7848e-39 = inf
	(b"11011000001000010011010100011101", b"00000000000000000000000000000000"),
	(b"10000000010111010010011111101110", b"11011000001000010011010100011101"), -- -7.08998e+14 + -8.55503e-39 = -7.08998e+14
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110111010111000110101", b"01111111100000000000000000000000"), -- inf + 5.48079e-39 = inf
	(b"11100010100110101110100000001111", b"00000000000000000000000000000000"),
	(b"00000000010101011101010110101011", b"11100010100110101110100000001111"), -- -1.42876e+21 + 7.88267e-39 = -1.42876e+21
	(b"01010111101110011110110011011000", b"00000000000000000000000000000000"),
	(b"00000000011101111010000000100110", b"01010111101110011110110011011000"), -- 4.08854e+14 + 1.09859e-38 = 4.08854e+14
	(b"01101000101101011111100001010010", b"00000000000000000000000000000000"),
	(b"10000000000011101011011001000011", b"01101000101101011111100001010010"), -- 6.87463e+24 + -1.35108e-39 = 6.87463e+24
	(b"01001101010001110010101100001100", b"00000000000000000000000000000000"),
	(b"00000000010111110011000111000101", b"01001101010001110010101100001100"), -- 2.08843e+08 + 8.74223e-39 = 2.08843e+08
	(b"01000000000101100011001110010100", b"00000000000000000000000000000000"),
	(b"10000000010010110001101011101110", b"01000000000101100011001110010100"), -- 2.3469 + -6.89732e-39 = 2.3469
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100100111000000100001", b"00000000000100100111000000100001"), -- 0 + 1.69326e-39 = 1.69326e-39
	(b"10011010100001000010101011111000", b"00000000000000000000000000000000"),
	(b"10000000010101010001111010110110", b"10011010100001000010101011111000"), -- -5.46633e-23 + -7.81703e-39 = -5.46633e-23
	(b"11000110011000001001110101111101", b"00000000000000000000000000000000"),
	(b"10000000011011000011001011010110", b"11000110011000001001110101111101"), -- -14375.4 + -9.93647e-39 = -14375.4
	(b"00011101101111111001100100110110", b"00000000000000000000000000000000"),
	(b"10000000001011000001010000110110", b"00011101101111111001100100110110"), -- 5.07157e-21 + -4.04801e-39 = 5.07157e-21
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111010001010001110010", b"00000000000111010001010001110010"), -- -0 + 2.67056e-39 = 2.67056e-39
	(b"11100001100110010010011011011111", b"00000000000000000000000000000000"),
	(b"10000000001001001111111000111000", b"11100001100110010010011011011111"), -- -3.53144e+20 + -3.39727e-39 = -3.53144e+20
	(b"11000111000011000000010001100011", b"00000000000000000000000000000000"),
	(b"00000000001011001111101100111001", b"11000111000011000000010001100011"), -- -35844.4 + 4.13088e-39 = -35844.4
	(b"10000000000000000000000100010011", b"00000000000000000000000000000000"),
	(b"00000000010111011111111100101111", b"00000000010111011111111000011100"), -- -3.85357e-43 + 8.63224e-39 = 8.63186e-39
	(b"11001010011011110001000000110110", b"00000000000000000000000000000000"),
	(b"00000000000011011011001101110010", b"11001010011011110001000000110110"), -- -3.91681e+06 + 1.25823e-39 = -3.91681e+06
	(b"11100011011011011101011111010100", b"00000000000000000000000000000000"),
	(b"00000000001101011010000100011101", b"11100011011011011101011111010100"), -- -4.38743e+21 + 4.92508e-39 = -4.38743e+21
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110101101101100000101", b"11111111100000000000000000000000"), -- -inf + 5.40503e-39 = -inf
	(b"11110111110001011110010110001110", b"00000000000000000000000000000000"),
	(b"00000000000010111101111110110111", b"11110111110001011110010110001110"), -- -8.02764e+33 + 1.09044e-39 = -8.02764e+33
	(b"01010110101111110110010110100111", b"00000000000000000000000000000000"),
	(b"00000000011010011110010111000010", b"01010110101111110110010110100111"), -- 1.05222e+14 + 9.72515e-39 = 1.05222e+14
	(b"11110000101111001110010000110110", b"00000000000000000000000000000000"),
	(b"10000000000110010101110011011010", b"11110000101111001110010000110110"), -- -4.67673e+29 + -2.3292e-39 = -4.67673e+29
	(b"01100001010101111100011100110001", b"00000000000000000000000000000000"),
	(b"00000000001000110011100000101100", b"01100001010101111100011100110001"), -- 2.48775e+20 + 3.23439e-39 = 2.48775e+20
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011110101111011111000", b"11111111100000000000000000000000"), -- -inf + 1.4116e-39 = -inf
	(b"01001011111110101011000111101110", b"00000000000000000000000000000000"),
	(b"10000000011001111000000010101111", b"01001011111110101011000111101110"), -- 3.28591e+07 + -9.50522e-39 = 3.28591e+07
	(b"10010101111110111100110010110001", b"00000000000000000000000000000000"),
	(b"10000000001101010110101010110001", b"10010101111110111100110010110001"), -- -1.01701e-25 + -4.90555e-39 = -1.01701e-25
	(b"00111111110101101000000100000110", b"00000000000000000000000000000000"),
	(b"00000000000110111100000011110011", b"00111111110101101000000100000110"), -- 1.67581 + 2.54878e-39 = 1.67581
	(b"00000011101000011000100011111111", b"00000000000000000000000000000000"),
	(b"00000000001000101110111101110011", b"00000011101000100001010010111101"), -- 9.49418e-37 + 3.20831e-39 = 9.52627e-37
	(b"01100010111100111001000110110110", b"00000000000000000000000000000000"),
	(b"10000000011110000111010110001001", b"01100010111100111001000110110110"), -- 2.24653e+21 + -1.10624e-38 = 2.24653e+21
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010010111001011101010110", b"10000000010010111001011101010110"), -- -0 + -6.94195e-39 = -6.94195e-39
	(b"10100000001000010111101100111001", b"00000000000000000000000000000000"),
	(b"00000000011111100000100101010101", b"10100000001000010111101100111001"), -- -1.3678e-19 + 1.15746e-38 = -1.3678e-19
	(b"01100000010101001100001100000111", b"00000000000000000000000000000000"),
	(b"10000000000000101110101100100101", b"01100000010101001100001100000111"), -- 6.13244e+19 + -2.68025e-40 = 6.13244e+19
	(b"10010100100000111011010001111110", b"00000000000000000000000000000000"),
	(b"00000000011011001110101010100111", b"10010100100000111011010001111110"), -- -1.32988e-26 + 1.00024e-38 = -1.32988e-26
	(b"11100101000110111101100110100100", b"00000000000000000000000000000000"),
	(b"00000000011110110110100110000110", b"11100101000110111101100110100100"), -- -4.59988e+22 + 1.13336e-38 = -4.59988e+22
	(b"11110111110100000100000011011011", b"00000000000000000000000000000000"),
	(b"00000000011000011100110111110010", b"11110111110100000100000011011011"), -- -8.44776e+33 + 8.98192e-39 = -8.44776e+33
	(b"11000101100011011000010110110010", b"00000000000000000000000000000000"),
	(b"10000000001100110010111000101101", b"11000101100011011000010110110010"), -- -4528.71 + -4.70018e-39 = -4528.71
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010000101111110010000101", b"01111111100000000000000000000000"), -- inf + 6.15173e-39 = inf
	(b"00111000011011001010011101000100", b"00000000000000000000000000000000"),
	(b"00000000000010111010110011010100", b"00111000011011001010011101000100"), -- 5.64226e-05 + 1.07219e-39 = 5.64226e-05
	(b"00000000000000000000000011010101", b"00000000000000000000000000000000"),
	(b"00000000001011001100101101101111", b"00000000001011001100110001000100"), -- 2.98477e-43 + 4.11374e-39 = 4.11404e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101001011100001000101", b"01111111100000000000000000000000"), -- inf + -4.84155e-39 = inf
	(b"11010101001111111100001001100001", b"00000000000000000000000000000000"),
	(b"10000000011110011101101000000000", b"11010101001111111100001001100001"), -- -1.31776e+13 + -1.11903e-38 = -1.31776e+13
	(b"00011100101110001011011101101000", b"00000000000000000000000000000000"),
	(b"10000000000001101000011000111111", b"00011100101110001011011101101000"), -- 1.22235e-21 + -5.99171e-40 = 1.22235e-21
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010010110101010101001101", b"10000000010010110101010101001101"), -- 0 + -6.91826e-39 = -6.91826e-39
	(b"00100010101000011110111101111000", b"00000000000000000000000000000000"),
	(b"00000000011001100100011001010110", b"00100010101000011110111101111000"), -- 4.38927e-18 + 9.39245e-39 = 4.38927e-18
	(b"00101111110110010101100111100001", b"00000000000000000000000000000000"),
	(b"10000000000011010011010000000000", b"00101111110110010101100111100001"), -- 3.95359e-10 + -1.21252e-39 = 3.95359e-10
	(b"11110001001011000101011000110110", b"00000000000000000000000000000000"),
	(b"00000000001001111101001110110000", b"11110001001011000101011000110110"), -- -8.5337e+29 + 3.65752e-39 = -8.5337e+29
	(b"10000000000000000000000000000101", b"00000000000000000000000000000000"),
	(b"10000000010010111010111010101111", b"10000000010010111010111010110100"), -- -7.00649e-45 + -6.95033e-39 = -6.95033e-39
	(b"00001110100001111110101000000001", b"00000000000000000000000000000000"),
	(b"00000000011100101111000000111010", b"00001110100001111110101000000001"), -- 3.35054e-30 + 1.05554e-38 = 3.35054e-30
	(b"01101001101010010111010000000011", b"00000000000000000000000000000000"),
	(b"10000000001000010111011011001111", b"01101001101010010111010000000011"), -- 2.5607e+25 + -3.07319e-39 = 2.5607e+25
	(b"00010110001100100110101010111001", b"00000000000000000000000000000000"),
	(b"00000000001000011010100011100001", b"00010110001100100110101010111001"), -- 1.44124e-25 + 3.09115e-39 = 1.44124e-25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110010100100110011010", b"11111111100000000000000000000000"), -- -inf + -5.26103e-39 = -inf
	(b"11010110111001100110000000011011", b"00000000000000000000000000000000"),
	(b"10000000011110101000101110110101", b"11010110111001100110000000011011"), -- -1.2665e+14 + -1.1254e-38 = -1.2665e+14
	(b"10001111011111001000111001111000", b"00000000000000000000000000000000"),
	(b"00000000010100010101100000001110", b"10001111011111001000111001111000"), -- -1.2452e-29 + 7.47026e-39 = -1.2452e-29
	(b"01110001000100110110100110111111", b"00000000000000000000000000000000"),
	(b"10000000001000001011100001001100", b"01110001000100110110100110111111"), -- 7.29954e+29 + -3.00485e-39 = 7.29954e+29
	(b"00110110010000100001101010001100", b"00000000000000000000000000000000"),
	(b"00000000011100101100111100010110", b"00110110010000100001101010001100"), -- 2.89237e-06 + 1.05435e-38 = 2.89237e-06
	(b"00011111001001111000100011111011", b"00000000000000000000000000000000"),
	(b"00000000000110011111000010101000", b"00011111001001111000100011111011"), -- 3.54769e-20 + 2.38222e-39 = 3.54769e-20
	(b"01000101000000010101011000100110", b"00000000000000000000000000000000"),
	(b"10000000010010000111110010101000", b"01000101000000010101011000100110"), -- 2069.38 + -6.65687e-39 = 2069.38
	(b"00010101001011110100101110111101", b"00000000000000000000000000000000"),
	(b"10000000010100100001100000101110", b"00010101001011110100101110111101"), -- 3.54007e-26 + -7.53918e-39 = 3.54007e-26
	(b"00100011000100101011010001001000", b"00000000000000000000000000000000"),
	(b"00000000011101110100010001100000", b"00100011000100101011010001001000"), -- 7.95285e-18 + 1.0953e-38 = 7.95285e-18
	(b"10110000001110011111010100011111", b"00000000000000000000000000000000"),
	(b"10000000000110100000110110111000", b"10110000001110011111010100011111"), -- -6.76509e-10 + -2.39264e-39 = -6.76509e-10
	(b"00110110001101000111000010001101", b"00000000000000000000000000000000"),
	(b"00000000000100101111100100010110", b"00110110001101000111000010001101"), -- 2.68876e-06 + 1.74239e-39 = 2.68876e-06
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011011011110001111110000", b"11111111100000000000000000000000"), -- -inf + -1.00918e-38 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010101001001110111101001", b"01111111100000000000000000000000"), -- inf + 7.77083e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010100111100100011001011", b"11111111100000000000000000000000"), -- -inf + 7.69438e-39 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001100100001100000111", b"00000000000001100100001100000111"), -- -0 + 5.75058e-40 = 5.75058e-40
	(b"11101001101010101111111111010001", b"00000000000000000000000000000000"),
	(b"10000000011100010111010011001100", b"11101001101010101111111111010001"), -- -2.58407e+25 + -1.04193e-38 = -2.58407e+25
	(b"11010111110000011111110001110010", b"00000000000000000000000000000000"),
	(b"00000000010111000101001001110101", b"11010111110000011111110001110010"), -- -4.2658e+14 + 8.47845e-39 = -4.2658e+14
	(b"11000101100001111100000011110100", b"00000000000000000000000000000000"),
	(b"00000000001100111101111101010110", b"11000101100001111100000011110100"), -- -4344.12 + 4.76373e-39 = -4344.12
	(b"11011110101110100000000110101111", b"00000000000000000000000000000000"),
	(b"10000000000001100111101110001100", b"11011110101110100000000110101111"), -- -6.70159e+18 + -5.95333e-40 = -6.70159e+18
	(b"10101110011011010100010101111101", b"00000000000000000000000000000000"),
	(b"10000000010001100100101001010011", b"10101110011011010100010101111101"), -- -5.39493e-11 + -6.45515e-39 = -5.39493e-11
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011111110010000100110010", b"00000000011111110010000100110010"), -- 0 + 1.1675e-38 = 1.1675e-38
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101110111000111000111", b"11111111100000000000000000000000"), -- -inf + 1.09692e-38 = -inf
	(b"00111111101011001001110010111010", b"00000000000000000000000000000000"),
	(b"10000000010100001011000110100110", b"00111111101011001001110010111010"), -- 1.34853 + -7.41057e-39 = 1.34853
	(b"00111101101000101100010001111011", b"00000000000000000000000000000000"),
	(b"10000000010010111100111101100000", b"00111101101000101100010001111011"), -- 0.0794763 + -6.96205e-39 = 0.0794763
	(b"00011110101010010111000010010001", b"00000000000000000000000000000000"),
	(b"00000000000100011100100001101110", b"00011110101010010111000010010001"), -- 1.79401e-20 + 1.6331e-39 = 1.79401e-20
	(b"10100110001101110010011011010100", b"00000000000000000000000000000000"),
	(b"10000000011100010100000101101111", b"10100110001101110010011011010100"), -- -6.35435e-16 + -1.04009e-38 = -6.35435e-16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110001101101100110010", b"01111111100000000000000000000000"), -- inf + -8.16016e-39 = inf
	(b"00100110011110000000111111011011", b"00000000000000000000000000000000"),
	(b"00000000011000100110010111100011", b"00100110011110000000111111011011"), -- 8.60638e-16 + 9.03643e-39 = 8.60638e-16
	(b"10000000000000101111001101111100", b"00000000000000000000000000000000"),
	(b"00000000010111100010101000110111", b"00000000010110110011011010111011"), -- -2.71017e-40 + 8.64768e-39 = 8.37666e-39
	(b"11011101101100011010010010011010", b"00000000000000000000000000000000"),
	(b"10000000011001101101101110011010", b"11011101101100011010010010011010"), -- -1.60007e+18 + -9.446e-39 = -1.60007e+18
	(b"10111001010000000111110011101010", b"00000000000000000000000000000000"),
	(b"00000000010000110011000100101111", b"10111001010000000111110011101010"), -- -0.000183571 + 6.17062e-39 = -0.000183571
	(b"00110000010010000100111111111000", b"00000000000000000000000000000000"),
	(b"00000000010101111000001010000011", b"00110000010010000100111111111000"), -- 7.28732e-10 + 8.03651e-39 = 7.28732e-10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011000101100101010001001", b"11111111100000000000000000000000"), -- -inf + 9.07253e-39 = -inf
	(b"10101110001001101010001001100011", b"00000000000000000000000000000000"),
	(b"10000000001101100011001111110101", b"10101110001001101010001001100011"), -- -3.78883e-11 + -4.97776e-39 = -3.78883e-11
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011010110001010011011101", b"10000000011010110001010011011101"), -- -0 + -9.83388e-39 = -9.83388e-39
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"00000000011110001000010001011001", b"00000000011110001000010001011000"), -- -1.4013e-45 + 1.10677e-38 = 1.10677e-38
	(b"01100110110011100101011110000011", b"00000000000000000000000000000000"),
	(b"00000000010001111101011100101000", b"01100110110011100101011110000011"), -- 4.87211e+23 + 6.5975e-39 = 4.87211e+23
	(b"00000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"00000000010100101110100101011010", b"00000000010100101110100101011011"), -- 1.4013e-45 + 7.61422e-39 = 7.61422e-39
	(b"11101101100001101100001111000111", b"00000000000000000000000000000000"),
	(b"00000000001011111111111111100111", b"11101101100001101100001111000111"), -- -5.21346e+27 + 4.40807e-39 = -5.21346e+27
	(b"00101110100110110110011001101010", b"00000000000000000000000000000000"),
	(b"10000000000010001010110000101000", b"00101110100110110110011001101010"), -- 7.06678e-11 + -7.96442e-40 = 7.06678e-11
	(b"00100100000000101111001111101001", b"00000000000000000000000000000000"),
	(b"00000000001110001011000100010110", b"00100100000000101111001111101001"), -- 2.83959e-17 + 5.20631e-39 = 2.83959e-17
	(b"00100111101101110011011001011111", b"00000000000000000000000000000000"),
	(b"00000000000111001110110110011101", b"00100111101101110011011001011111"), -- 5.08517e-15 + 2.65663e-39 = 5.08517e-15
	(b"10111100011110111001010011110000", b"00000000000000000000000000000000"),
	(b"00000000011001101100001000001100", b"10111100011110111001010011110000"), -- -0.0153553 + 9.43683e-39 = -0.0153553
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111010000101011100100", b"11111111100000000000000000000000"), -- -inf + 5.60587e-39 = -inf
	(b"00010011111100000100011011010000", b"00000000000000000000000000000000"),
	(b"00000000010011101000001000110011", b"00010011111100000100011011010000"), -- 6.06543e-27 + 7.20988e-39 = 6.06543e-27
	(b"01000100010110101100101000001001", b"00000000000000000000000000000000"),
	(b"10000000000011001110010110110101", b"01000100010110101100101000001001"), -- 875.157 + -1.18443e-39 = 875.157
	(b"11101111001001010100011010100110", b"00000000000000000000000000000000"),
	(b"00000000001001110100110110110101", b"11101111001001010100011010100110"), -- -5.11504e+28 + 3.60946e-39 = -5.11504e+28
	(b"10000101101110011100100000010011", b"00000000000000000000000000000000"),
	(b"00000000011101100000101001011011", b"10000101101110011010101010010000"), -- -1.74708e-35 + 1.08403e-38 = -1.746e-35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010010000110111000100000", b"11111111100000000000000000000000"), -- -inf + 6.65166e-39 = -inf
	(b"00101110111111101100001111111011", b"00000000000000000000000000000000"),
	(b"10000000001111010011110101101001", b"00101110111111101100001111111011"), -- 1.15854e-10 + -5.624e-39 = 1.15854e-10
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010000110000101100000011", b"00000000010000110000101100000011"), -- -0 + 6.15693e-39 = 6.15693e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001101101111111101010001", b"00000000001101101111111101010001"), -- -0 + 5.05071e-39 = 5.05071e-39
	(b"11000111000011011100101000111010", b"00000000000000000000000000000000"),
	(b"00000000010111010111010111000111", b"11000111000011011100101000111010"), -- -36298.2 + 8.58295e-39 = -36298.2
	(b"01000111111100110101111010110100", b"00000000000000000000000000000000"),
	(b"10000000000010001101001011000101", b"01000111111100110101111010110100"), -- 124605 + -8.10294e-40 = 124605
	(b"00100011111100000011110011110111", b"00000000000000000000000000000000"),
	(b"10000000001100100001110010111011", b"00100011111100000011110011110111"), -- 2.60467e-17 + -4.60208e-39 = 2.60467e-17
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010001110100010010000", b"00000000000010001110100010010000"), -- 0 + 8.18112e-40 = 8.18112e-40
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101110100100111001111", b"11111111100000000000000000000000"), -- -inf + -1.09549e-38 = -inf
	(b"01001111110001010000111111110111", b"00000000000000000000000000000000"),
	(b"00000000001101001111100010011000", b"01001111110001010000111111110111"), -- 6.61232e+09 + 4.86462e-39 = 6.61232e+09
	(b"11000100101101000100110110011100", b"00000000000000000000000000000000"),
	(b"10000000011101101010111111001100", b"11000100101101000100110110011100"), -- -1442.43 + -1.08997e-38 = -1442.43
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011111010001000011011110", b"11111111100000000000000000000000"), -- -inf + -1.14855e-38 = -inf
	(b"10101011000110001011011110000001", b"00000000000000000000000000000000"),
	(b"10000000001110010011011011111110", b"10101011000110001011011110000001"), -- -5.42559e-13 + -5.25435e-39 = -5.42559e-13
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000111111011100111110", b"10000000011000111111011100111110"), -- -0 + -9.18041e-39 = -9.18041e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100000000001110001110", b"00000000000100000000001110001110"), -- -0 + 1.47064e-39 = 1.47064e-39
	(b"10100000001011110111001100010110", b"00000000000000000000000000000000"),
	(b"10000000011110001101011110111011", b"10100000001011110111001100010110"), -- -1.48612e-19 + -1.10976e-38 = -1.48612e-19
	(b"01010001101100110000111100111001", b"00000000000000000000000000000000"),
	(b"00000000000001010001010111110100", b"01010001101100110000111100111001"), -- 9.61318e+10 + 4.67053e-40 = 9.61318e+10
	(b"11110011010101010101100111010011", b"00000000000000000000000000000000"),
	(b"00000000010110010011100010101011", b"11110011010101010101100111010011"), -- -1.69034e+31 + 8.19369e-39 = -1.69034e+31
	(b"11010111010001101101100110000101", b"00000000000000000000000000000000"),
	(b"10000000001111111010101111010011", b"11010111010001101101100110000101"), -- -2.18638e+14 + -5.84728e-39 = -2.18638e+14
	(b"10010111100000011000011110110001", b"00000000000000000000000000000000"),
	(b"10000000000000010010011001010001", b"10010111100000011000011110110001"), -- -8.37068e-25 + -1.05581e-40 = -8.37068e-25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011001110110001101000", b"11111111100000000000000000000000"), -- -inf + 1.0003e-38 = -inf
	(b"10010000001111100011010110000111", b"00000000000000000000000000000000"),
	(b"10000000010111011000001000101111", b"10010000001111100011010110000111"), -- -3.75121e-29 + -8.5874e-39 = -3.75121e-29
	(b"11101011100010001011111010001000", b"00000000000000000000000000000000"),
	(b"00000000000101111010101110000110", b"11101011100010001011111010001000"), -- -3.30627e+26 + 2.17375e-39 = -3.30627e+26
	(b"10000000000000000000000101110010", b"00000000000000000000000000000000"),
	(b"10000000000101101000111001111101", b"10000000000101101000111111101111"), -- -5.1848e-43 + -2.0715e-39 = -2.07201e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010011111100010100111101", b"11111111100000000000000000000000"), -- -inf + 7.32576e-39 = -inf
	(b"00001011000011101100000011101111", b"00000000000000000000000000000000"),
	(b"10000000010000000101101000101111", b"00001011000011101100000011101101"), -- 2.74934e-32 + -5.90982e-39 = 2.74933e-32
	(b"00111100101011010010011010111110", b"00000000000000000000000000000000"),
	(b"00000000001100010110110100101110", b"00111100101011010010011010111110"), -- 0.0211366 + 4.53911e-39 = 0.0211366
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111100101110001001100", b"01111111100000000000000000000000"), -- inf + -8.66565e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000010000010100000111", b"00000000001000010000010100000111"), -- 0 + 3.03237e-39 = 3.03237e-39
	(b"00010111101100101010100101001011", b"00000000000000000000000000000000"),
	(b"00000000000100000101110111100100", b"00010111101100101010100101001011"), -- 1.15457e-24 + 1.50305e-39 = 1.15457e-24
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011001000111100110010", b"00000000001011001000111100110010"), -- 0 + 4.09213e-39 = 4.09213e-39
	(b"01000110011100110101011110111001", b"00000000000000000000000000000000"),
	(b"10000000000001001000011111011101", b"01000110011100110101011110111001"), -- 15573.9 + -4.16081e-40 = 15573.9
	(b"10100001000001000011110101010001", b"00000000000000000000000000000000"),
	(b"00000000011010010011111110010010", b"10100001000001000011110101010001"), -- -4.48045e-19 + 9.66553e-39 = -4.48045e-19
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100010111111111000010", b"00000000000100010111111111000010"), -- -0 + 1.60703e-39 = 1.60703e-39
	(b"00111111111111101011011100011011", b"00000000000000000000000000000000"),
	(b"00000000001010110100101101101111", b"00111111111111101011011100011011"), -- 1.98996 + 3.97599e-39 = 1.98996
	(b"11111000001001001010011001100110", b"00000000000000000000000000000000"),
	(b"00000000001010110001010100001011", b"11111000001001001010011001100110"), -- -1.3358e+34 + 3.95648e-39 = -1.3358e+34
	(b"00011011101000001111011000111110", b"00000000000000000000000000000000"),
	(b"00000000010111010000111101101111", b"00011011101000001111011000111110"), -- 2.66289e-22 + 8.54624e-39 = 2.66289e-22
	(b"10101010011101000100010100100111", b"00000000000000000000000000000000"),
	(b"00000000000110000001110100110011", b"10101010011101000100010100100111"), -- -2.16955e-13 + 2.21453e-39 = -2.16955e-13
	(b"10001001110101111000110000100000", b"00000000000000000000000000000000"),
	(b"00000000010000110011101100000010", b"10001001110101111000110000001111"), -- -5.18911e-33 + 6.17415e-39 = -5.18911e-33
	(b"01001100000110101011010010001111", b"00000000000000000000000000000000"),
	(b"00000000011010101111101011011001", b"01001100000110101011010010001111"), -- 4.05551e+07 + 9.82455e-39 = 4.05551e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001111110111111101010", b"00000000011001111110111111101010"), -- -0 + 9.54512e-39 = 9.54512e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100100010111111100101", b"11111111100000000000000000000000"), -- -inf + -1.04864e-38 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011110110000011001001101", b"11111111100000000000000000000000"), -- -inf + 1.1298e-38 = -inf
	(b"11110110100111101010011111111110", b"00000000000000000000000000000000"),
	(b"10000000000010101010100111000101", b"11110110100111101010011111111110"), -- -1.60897e+33 + -9.79257e-40 = -1.60897e+33
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010000011001000001010000", b"11111111100000000000000000000000"), -- -inf + 6.02108e-39 = -inf
	(b"10111110001011011101000101110101", b"00000000000000000000000000000000"),
	(b"00000000010001111010011001011111", b"10111110001011011101000101110101"), -- -0.169744 + 6.58e-39 = -0.169744
	(b"10101011111101011001000110110100", b"00000000000000000000000000000000"),
	(b"10000000011001110101111111011110", b"10101011111101011001000110110100"), -- -1.74487e-12 + -9.49345e-39 = -1.74487e-12
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000001100100111111101", b"10000000011000001100100111111101"), -- 0 + -8.88867e-39 = -8.88867e-39
	(b"10101011010010001111011001011110", b"00000000000000000000000000000000"),
	(b"00000000001000100000000001011110", b"10101011010010001111011001011110"), -- -7.13962e-13 + 3.12254e-39 = -7.13962e-13
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001100101101111101000100", b"00000000001100101101111101000100"), -- 0 + 4.67187e-39 = 4.67187e-39
	(b"11101000110101001111101001110100", b"00000000000000000000000000000000"),
	(b"10000000001010011011000110000001", b"11101000110101001111101001110100"), -- -8.04609e+24 + -3.82893e-39 = -8.04609e+24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010011001010101011001101", b"00000000010011001010101011001101"), -- -0 + 7.04077e-39 = 7.04077e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011111101110110100000101", b"11111111100000000000000000000000"), -- -inf + -1.16563e-38 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001001010011000001110", b"11111111100000000000000000000000"), -- -inf + -9.24312e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110010010101000000010", b"01111111100000000000000000000000"), -- inf + -5.24969e-39 = inf
	(b"11110000000110010100100101110101", b"00000000000000000000000000000000"),
	(b"00000000000100111111101110001000", b"11110000000110010100100101110101"), -- -1.8976e+29 + 1.83511e-39 = -1.8976e+29
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011111011010011000110", b"01111111100000000000000000000000"), -- inf + 1.44238e-39 = inf
	(b"01011111101111100011101001110001", b"00000000000000000000000000000000"),
	(b"00000000011011101100101001100011", b"01011111101111100011101001110001"), -- 2.74148e+19 + 1.01745e-38 = 2.74148e+19
	(b"01010110101100101011000011000100", b"00000000000000000000000000000000"),
	(b"10000000010000000100101100100001", b"01010110101100101011000011000100"), -- 9.82361e+13 + -5.90442e-39 = 9.82361e+13
	(b"11010010101111011001001000000001", b"00000000000000000000000000000000"),
	(b"00000000001111011000111110011011", b"11010010101111011001001000000001"), -- -4.07099e+11 + 5.65348e-39 = -4.07099e+11
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010011101001110111101000", b"00000000010011101001110111101000"), -- 0 + 7.21981e-39 = 7.21981e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111101001110101001100", b"01111111100000000000000000000000"), -- inf + 5.75023e-39 = inf
	(b"00000000000000001010110111101101", b"00000000000000000000000000000000"),
	(b"10000000011111100110111110010111", b"10000000011111011100000110101010"), -- 6.23928e-41 + -1.16113e-38 = -1.15489e-38
	(b"11011101001110110000111111011010", b"00000000000000000000000000000000"),
	(b"00000000010000110100011000010101", b"11011101001110110000111111011010"), -- -8.42452e+17 + 6.17812e-39 = -8.42452e+17
	(b"00000000110010001010100101011101", b"00000000000000000000000000000000"),
	(b"00000000010110111111100001100100", b"00000001000100100101000011100000"), -- 1.84279e-38 + 8.44614e-39 = 2.6874e-38
	(b"01000110101011101110011100000010", b"00000000000000000000000000000000"),
	(b"00000000001111010000000011000110", b"01000110101011101110011100000010"), -- 22387.5 + 5.60224e-39 = 22387.5
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111010011110000000101", b"11111111100000000000000000000000"), -- -inf + 5.6235e-39 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010000100010101110010", b"00000000000010000100010101110010"), -- -0 + 7.59596e-40 = 7.59596e-40
	(b"00000000000000000000000000010011", b"00000000000000000000000000000000"),
	(b"00000000000101100110110001100010", b"00000000000101100110110001110101"), -- 2.66247e-44 + 2.05926e-39 = 2.05929e-39
	(b"01101111010100101001100011111010", b"00000000000000000000000000000000"),
	(b"00000000010110101001101011010000", b"01101111010100101001100011111010"), -- 6.51768e+28 + 8.32073e-39 = 6.51768e+28
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010100111000011011011", b"11111111100000000000000000000000"), -- -inf + -3.89758e-39 = -inf
	(b"00100110101010110001101000010011", b"00000000000000000000000000000000"),
	(b"10000000011000001101010111100000", b"00100110101010110001101000010011"), -- 1.18726e-15 + -8.89293e-39 = 1.18726e-15
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010100001100100011110010", b"01111111100000000000000000000000"), -- inf + -7.41893e-39 = inf
	(b"10110100010001110100100110001010", b"00000000000000000000000000000000"),
	(b"00000000001001110000011110100011", b"10110100010001110100100110001010"), -- -1.85601e-07 + 3.58432e-39 = -1.85601e-07
	(b"00000000000110100100100001111100", b"00000000000000000000000000000000"),
	(b"10000000011010111010000000010010", b"10000000010100010101011110010110"), -- 2.41373e-39 + -9.88382e-39 = -7.4701e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101000000100111110100", b"11111111100000000000000000000000"), -- -inf + 1.06565e-38 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000001101101101100010100", b"10000000000001101101101100010100"), -- -0 + -6.29603e-40 = -6.29603e-40
	(b"10101111010000100111001100001101", b"00000000000000000000000000000000"),
	(b"10000000010101111010111111100010", b"10101111010000100111001100001101"), -- -1.76851e-10 + -8.05278e-39 = -1.76851e-10
	(b"01010111100000100110101100101000", b"00000000000000000000000000000000"),
	(b"10000000000001000000011000101111", b"01010111100000100110101100101000"), -- 2.86793e+14 + -3.6956e-40 = 2.86793e+14
	(b"11001000111100001111110000000001", b"00000000000000000000000000000000"),
	(b"00000000011100010011101001001111", b"11001000111100001111110000000001"), -- -493536 + 1.03983e-38 = -493536
	(b"01110001101011011011110101100111", b"00000000000000000000000000000000"),
	(b"00000000001101110110100111001110", b"01110001101011011011110101100111"), -- 1.72064e+30 + 5.08891e-39 = 1.72064e+30
	(b"11110110110110010110111100010010", b"00000000000000000000000000000000"),
	(b"10000000010010010000111101101001", b"11110110110110010110111100010010"), -- -2.20504e+33 + -6.70952e-39 = -2.20504e+33
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111011000111010001010", b"00000000000111011000111010001010"), -- 0 + 2.71436e-39 = 2.71436e-39
	(b"01000100011011111011111110111011", b"00000000000000000000000000000000"),
	(b"10000000000001100111110100000100", b"01000100011011111011111110111011"), -- 958.996 + -5.9586e-40 = 958.996
	(b"10001100001101001100011110001010", b"00000000000000000000000000000000"),
	(b"00000000000111001100011011101111", b"10001100001101001100011110001010"), -- -1.39267e-31 + 2.64276e-39 = -1.39267e-31
	(b"01110101100111001100010011010000", b"00000000000000000000000000000000"),
	(b"10000000011100100001000100011111", b"01110101100111001100010011010000"), -- 3.97456e+32 + -1.04754e-38 = 3.97456e+32
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100111010111110100000", b"01111111100000000000000000000000"), -- inf + 1.80788e-39 = inf
	(b"10001011101110111001010110010101", b"00000000000000000000000000000000"),
	(b"10000000000110101001011011011010", b"10001011101110111001010110010101"), -- -7.22548e-32 + -2.44184e-39 = -7.22548e-32
	(b"00000000000000000000000000101001", b"00000000000000000000000000000000"),
	(b"10000000001001000111101101000010", b"10000000001001000111101100011001"), -- 5.74532e-44 + -3.35029e-39 = -3.35024e-39
	(b"00111110100100100000011100001100", b"00000000000000000000000000000000"),
	(b"00000000011011101010000001000011", b"00111110100100100000011100001100"), -- 0.28521 + 1.01594e-38 = 0.28521
	(b"11111001011100011101010101011001", b"00000000000000000000000000000000"),
	(b"00000000001001011101011000011010", b"11111001011100011101010101011001"), -- -7.84794e+34 + 3.47472e-39 = -7.84794e+34
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000101000010000001011111", b"01111111100000000000000000000000"), -- inf + 1.84832e-39 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001010111110001000001", b"00000000011001010111110001000001"), -- -0 + 9.31996e-39 = 9.31996e-39
	(b"11100100100111100011010001111111", b"00000000000000000000000000000000"),
	(b"00000000001010111010110101111100", b"11100100100111100011010001111111"), -- -2.33469e+22 + 4.01116e-39 = -2.33469e+22
	(b"11111010001101100100011100010111", b"00000000000000000000000000000000"),
	(b"10000000010011110010010000100011", b"11111010001101100100011100010111"), -- -2.3661e+35 + -7.26797e-39 = -2.3661e+35
	(b"01010100111101000010111110111010", b"00000000000000000000000000000000"),
	(b"00000000001111110111010001110111", b"01010100111101000010111110111010"), -- 8.39018e+12 + 5.82742e-39 = 8.39018e+12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001100100010110111010000", b"11111111100000000000000000000000"), -- -inf + 4.60821e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101010011100011011010", b"11111111100000000000000000000000"), -- -inf + -4.88768e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010101100001111101100", b"01111111100000000000000000000000"), -- inf + -3.92737e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000011110001111110010", b"01111111100000000000000000000000"), -- inf + 1.73607e-40 = inf
	(b"01100011000100110110001111000101", b"00000000000000000000000000000000"),
	(b"10000000001010100011010101000110", b"01100011000100110110001111000101"), -- 2.71886e+21 + -3.8762e-39 = 2.71886e+21
	(b"01010110001100101000001011110110", b"00000000000000000000000000000000"),
	(b"10000000001011100111001111010001", b"01010110001100101000001011110110"), -- 4.90689e+13 + -4.26598e-39 = 4.90689e+13
	(b"10111110111001111111111101011010", b"00000000000000000000000000000000"),
	(b"10000000000000110000101100011110", b"10111110111001111111111101011010"), -- -0.45312 + -2.79495e-40 = -0.45312
	(b"11010100000010111011011101010010", b"00000000000000000000000000000000"),
	(b"10000000011100100001001110000110", b"11010100000010111011011101010010"), -- -2.4003e+12 + -1.04763e-38 = -2.4003e+12
	(b"01000010100001101101000001011100", b"00000000000000000000000000000000"),
	(b"00000000011011110111010000110001", b"01000010100001101101000001011100"), -- 67.407 + 1.02354e-38 = 67.407
	(b"01111011100101001111001011001010", b"00000000000000000000000000000000"),
	(b"00000000000111001011110101010000", b"01111011100101001111001011001010"), -- 1.54677e+36 + 2.63931e-39 = 1.54677e+36
	(b"11110000101000111001001101010010", b"00000000000000000000000000000000"),
	(b"10000000000011000011110000011000", b"11110000101000111001001101010010"), -- -4.04993e+29 + -1.12358e-39 = -4.04993e+29
	(b"11110111001011011101011100101110", b"00000000000000000000000000000000"),
	(b"10000000000110000101010000001101", b"11110111001011011101011100101110"), -- -3.52591e+33 + -2.2342e-39 = -3.52591e+33
	(b"11110010110001010001100101110100", b"00000000000000000000000000000000"),
	(b"10000000000111110100011001110100", b"11110010110001010001100101110100"), -- -7.80791e+30 + -2.87217e-39 = -7.80791e+30
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010010011101111101000100", b"10000000010010011101111101000100"), -- -0 + -6.78408e-39 = -6.78408e-39
	(b"00010111111101110010111010110000", b"00000000000000000000000000000000"),
	(b"10000000001010110000101011101001", b"00010111111101110010111010110000"), -- 1.59738e-24 + -3.95284e-39 = 1.59738e-24
	(b"11001100010100111100000000111011", b"00000000000000000000000000000000"),
	(b"10000000011101000100111001101011", b"11001100010100111100000000111011"), -- -5.55092e+07 + -1.0681e-38 = -5.55092e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110111001011000000011", b"00000000010110111001011000000011"), -- 0 + 8.41084e-39 = 8.41084e-39
	(b"10010000000100010110001101110000", b"00000000000000000000000000000000"),
	(b"10000000001001101111010010101101", b"10010000000100010110001101110000"), -- -2.86728e-29 + -3.57752e-39 = -2.86728e-29
	(b"11111011010001100101111000101100", b"00000000000000000000000000000000"),
	(b"10000000010010000101010101010011", b"11111011010001100101111000101100"), -- -1.02998e+36 + -6.64276e-39 = -1.02998e+36
	(b"00010111000100110001100010001110", b"00000000000000000000000000000000"),
	(b"10000000011101000010010101011011", b"00010111000100110001100010001110"), -- 4.75293e-25 + -1.06663e-38 = 4.75293e-25
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100001001111010111010", b"01111111100000000000000000000000"), -- inf + -1.52631e-39 = inf
	(b"10101110110101000010111101001111", b"00000000000000000000000000000000"),
	(b"10000000010111010100000000000001", b"10101110110101000010111101001111"), -- -9.64905e-11 + -8.56366e-39 = -9.64905e-11
	(b"01011010100010000110001001111001", b"00000000000000000000000000000000"),
	(b"10000000000000010110111000100011", b"01011010100010000110001001111001"), -- 1.91944e+16 + -1.31345e-40 = 1.91944e+16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010111101001001011010", b"01111111100000000000000000000000"), -- inf + -1.08565e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001000010011110100010", b"10000000011001000010011110100010"), -- 0 + -9.19777e-39 = -9.19777e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001000011101110011111", b"10000000001001000011101110011111"), -- 0 + -3.32747e-39 = -3.32747e-39
	(b"00100110110010111000000110101011", b"00000000000000000000000000000000"),
	(b"00000000001100111000001001010100", b"00100110110010111000000110101011"), -- 1.41211e-15 + 4.73036e-39 = 1.41211e-15
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100110010101010110110", b"11111111100000000000000000000000"), -- -inf + -1.05764e-38 = -inf
	(b"11011010111111111011110100100010", b"00000000000000000000000000000000"),
	(b"00000000011100001000001001111110", b"11011010111111111011110100100010"), -- -3.5992e+16 + 1.03324e-38 = -3.5992e+16
	(b"11100110111000010110010111011101", b"00000000000000000000000000000000"),
	(b"00000000001111111111001011111011", b"11100110111000010110010111011101"), -- -5.32206e+23 + 5.8728e-39 = -5.32206e+23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010000011111010000001001", b"10000000010000011111010000001001"), -- 0 + -6.05685e-39 = -6.05685e-39
	(b"01010101101100110011010000111001", b"00000000000000000000000000000000"),
	(b"10000000010101101001100010110011", b"01010101101100110011010000111001"), -- 2.46296e+13 + -7.95263e-39 = 2.46296e+13
	(b"00010100001110111111101000000010", b"00000000000000000000000000000000"),
	(b"00000000000110000000100111100100", b"00010100001110111111101000000010"), -- 9.49039e-27 + 2.2076e-39 = 9.49039e-27
	(b"01100100001001000101110000101101", b"00000000000000000000000000000000"),
	(b"00000000000100000011010000100010", b"01100100001001000101110000101101"), -- 1.21276e+22 + 1.48807e-39 = 1.21276e+22
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110011110111100110110", b"11111111100000000000000000000000"), -- -inf + -1.11979e-38 = -inf
	(b"00101110011100110100100111111111", b"00000000000000000000000000000000"),
	(b"10000000010001101001001000100100", b"00101110011100110100100111111111"), -- 5.53175e-11 + -6.48091e-39 = 5.53175e-11
	(b"00001001100010001111100101000010", b"00000000000000000000000000000000"),
	(b"10000000000111000100010001010110", b"00001001100010001111100100111011"), -- 3.29752e-33 + -2.59591e-39 = 3.29752e-33
	(b"11011010010100111101111110101101", b"00000000000000000000000000000000"),
	(b"00000000000110010001010001101000", b"11011010010100111101111110101101"), -- -1.49093e+16 + 2.30321e-39 = -1.49093e+16
	(b"10000001001101000000011110001101", b"00000000000000000000000000000000"),
	(b"10000000000101100101110110111100", b"10000001001111110011011001101011"), -- -3.30662e-38 + -2.05401e-39 = -3.51202e-38
	(b"00110000001111010011111101100011", b"00000000000000000000000000000000"),
	(b"00000000000000000101110110101000", b"00110000001111010011111101100011"), -- 6.88479e-10 + 3.35975e-41 = 6.88479e-10
	(b"10101000000111100001000110100100", b"00000000000000000000000000000000"),
	(b"00000000010111010010100011110001", b"10101000000111100001000110100100"), -- -8.77459e-15 + 8.55539e-39 = -8.77459e-15
	(b"01110111010001100001110000101000", b"00000000000000000000000000000000"),
	(b"10000000011001001010001111011100", b"01110111010001100001110000101000"), -- 4.01815e+33 + -9.24233e-39 = 4.01815e+33
	(b"10001110101101000010111111111100", b"00000000000000000000000000000000"),
	(b"10000000010000001101001010000101", b"10001110101101000010111111111100"), -- -4.44196e-30 + -5.95299e-39 = -4.44196e-30
	(b"11101110101100010111101101100001", b"00000000000000000000000000000000"),
	(b"10000000001101011010110100010000", b"11101110101100010111101101100001"), -- -2.7464e+28 + -4.92936e-39 = -2.7464e+28
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010001101000000000011010", b"10000000010001101000000000011010"), -- -0 + -6.47444e-39 = -6.47444e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100010111111110100011", b"10000000011100010111111110100011"), -- -0 + -1.04232e-38 = -1.04232e-38
	(b"00111100111010110101110001010110", b"00000000000000000000000000000000"),
	(b"00000000000110011111011100001001", b"00111100111010110101110001010110"), -- 0.0287306 + 2.38451e-39 = 0.0287306
	(b"10110111000001111010011001100110", b"00000000000000000000000000000000"),
	(b"00000000001100100110111001110101", b"10110111000001111010011001100110"), -- -8.08537e-06 + 4.6314e-39 = -8.08537e-06
	(b"00000011111000001010000101110011", b"00000000000000000000000000000000"),
	(b"00000000000010100000010111110110", b"00000011111000001100100110001011"), -- 1.32026e-36 + 9.20493e-40 = 1.32118e-36
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011111100110101001000010", b"11111111100000000000000000000000"), -- -inf + -1.16094e-38 = -inf
	(b"10010100100101100010001000100000", b"00000000000000000000000000000000"),
	(b"00000000011001000010000100000111", b"10010100100101100010001000100000"), -- -1.51596e-26 + 9.1954e-39 = -1.51596e-26
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011111101110001001010111", b"11111111100000000000000000000000"), -- -inf + 1.16525e-38 = -inf
	(b"01101101010001100100111110001100", b"00000000000000000000000000000000"),
	(b"00000000011100110110010001101000", b"01101101010001100100111110001100"), -- 3.83589e+27 + 1.05971e-38 = 3.83589e+27
	(b"10100010011000010001101001000011", b"00000000000000000000000000000000"),
	(b"10000000010011010001111100010100", b"10100010011000010001101001000011"), -- -3.05071e-18 + -7.08248e-39 = -3.05071e-18
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010100101000101011111010", b"01111111100000000000000000000000"), -- inf + -7.58037e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100110100000111101000", b"11111111100000000000000000000000"), -- -inf + -1.76852e-39 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000001010101111000010100", b"10000000000001010101111000010100"), -- -0 + -4.92926e-40 = -4.92926e-40
	(b"11110110000011101000011111001101", b"00000000000000000000000000000000"),
	(b"00000000010100111111011001010010", b"11110110000011101000011111001101"), -- -7.22715e+32 + 7.71071e-39 = -7.22715e+32
	(b"00010001111111111101000011001001", b"00000000000000000000000000000000"),
	(b"00000000000000001100100001000101", b"00010001111111111101000011001001"), -- 4.03606e-28 + 7.18432e-41 = 4.03606e-28
	(b"00011011001101010111000000001101", b"00000000000000000000000000000000"),
	(b"10000000000000111000010111100110", b"00011011001101010111000000001101"), -- 1.50082e-22 + -3.2354e-40 = 1.50082e-22
	(b"10011000001001110011101000010010", b"00000000000000000000000000000000"),
	(b"10000000011001100000110111100001", b"10011000001001110011101000010010"), -- -2.16136e-24 + -9.3722e-39 = -2.16136e-24
	(b"01011010100100100110110100010000", b"00000000000000000000000000000000"),
	(b"00000000011000111011000011111100", b"01011010100100100110110100010000"), -- 2.06076e+16 + 9.1552e-39 = 2.06076e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100100001101000110001", b"11111111100000000000000000000000"), -- -inf + -1.66243e-39 = -inf
	(b"01110000100111111101000110110101", b"00000000000000000000000000000000"),
	(b"10000000001111001110100100001010", b"01110000100111111101000110110101"), -- 3.95693e+29 + -5.59373e-39 = 3.95693e+29
	(b"10100100000110110001010011111100", b"00000000000000000000000000000000"),
	(b"10000000001000011011001000010101", b"10100100000110110001010011111100"), -- -3.3628e-17 + -3.09446e-39 = -3.3628e-17
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010000010111001001010", b"01111111100000000000000000000000"), -- inf + -3.69003e-39 = inf
	(b"11011101001011000110111011110100", b"00000000000000000000000000000000"),
	(b"00000000010000100110111000111110", b"11011101001011000110111011110100"), -- -7.76571e+17 + 6.10069e-39 = -7.76571e+17
	(b"01011100101000011101001110010011", b"00000000000000000000000000000000"),
	(b"10000000001110100101010000111010", b"01011100101000011101001110010011"), -- 3.64401e+17 + -5.35667e-39 = 3.64401e+17
	(b"01100001110000000101101010000011", b"00000000000000000000000000000000"),
	(b"00000000011111100111000010111110", b"01100001110000000101101010000011"), -- 4.43537e+20 + 1.16117e-38 = 4.43537e+20
	(b"01010010000010101000000111011010", b"00000000000000000000000000000000"),
	(b"00000000011111100110101111001100", b"01010010000010101000000111011010"), -- 1.48721e+11 + 1.16099e-38 = 1.48721e+11
	(b"10011101100111011101011111000111", b"00000000000000000000000000000000"),
	(b"10000000000111110100100101010110", b"10011101100111011101011111000111"), -- -4.17807e-21 + -2.87321e-39 = -4.17807e-21
	(b"00101000101100111100011110101100", b"00000000000000000000000000000000"),
	(b"00000000011100110101101110101011", b"00101000101100111100011110101100"), -- 1.99596e-14 + 1.0594e-38 = 1.99596e-14
	(b"10000001001100011110000101101001", b"00000000000000000000000000000000"),
	(b"00000000001010111101110100000110", b"10000001000110111111001011100110"), -- -3.26715e-38 + 4.02821e-39 = -2.86433e-38
	(b"01101010000100000101000111001101", b"00000000000000000000000000000000"),
	(b"10000000010110101000010100010000", b"01101010000100000101000111001101"), -- 4.36179e+25 + -8.31293e-39 = 4.36179e+25
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011110010100011101001", b"00000000011011110010100011101001"), -- -0 + 1.02084e-38 = 1.02084e-38
	(b"11010011000001110001111100010101", b"00000000000000000000000000000000"),
	(b"00000000000100101111001011111011", b"11010011000001110001111100010101"), -- -5.80342e+11 + 1.7402e-39 = -5.80342e+11
	(b"10100010000000011111100101111111", b"00000000000000000000000000000000"),
	(b"00000000011110001000010001111001", b"10100010000000011111100101111111"), -- -1.76148e-18 + 1.10678e-38 = -1.76148e-18
	(b"11010000110110110100110110011000", b"00000000000000000000000000000000"),
	(b"10000000011101101110100100000001", b"11010000110110110100110110011000"), -- -2.94344e+10 + -1.09202e-38 = -2.94344e+10
	(b"00011010101001010010101011110001", b"00000000000000000000000000000000"),
	(b"10000000010001001110101100110101", b"00011010101001010010101011110001"), -- 6.83118e-23 + -6.32919e-39 = 6.83118e-23
	(b"01010011000010000011010101001101", b"00000000000000000000000000000000"),
	(b"00000000000100111110010000100010", b"01010011000010000011010101001101"), -- 5.8501e+11 + 1.82671e-39 = 5.8501e+11
	(b"11010000011001011000110100010111", b"00000000000000000000000000000000"),
	(b"00000000001000011110100110100011", b"11010000011001011000110100010111"), -- -1.54049e+10 + 3.11438e-39 = -1.54049e+10
	(b"00110000100011100011101001101111", b"00000000000000000000000000000000"),
	(b"00000000010110011000100100101011", b"00110000100011100011101001101111"), -- 1.03485e-09 + 8.22257e-39 = 1.03485e-09
	(b"11011011010110001111011100100101", b"00000000000000000000000000000000"),
	(b"10000000001001101101011111110100", b"11011011010110001111011100100101"), -- -6.10703e+16 + -3.56722e-39 = -6.10703e+16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011010011111000011011000", b"10000000011010011111000011011000"), -- 0 + -9.72913e-39 = -9.72913e-39
	(b"11011101101010011010000001100010", b"00000000000000000000000000000000"),
	(b"10000000010100001000110001100111", b"11011101101010011010000001100010"), -- -1.52786e+18 + -7.39721e-39 = -1.52786e+18
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011011110100011101001101", b"10000000011011110100011101001101"), -- 0 + -1.02193e-38 = -1.02193e-38
	(b"00111100100101101101011101100011", b"00000000000000000000000000000000"),
	(b"00000000010001101101000000011100", b"00111100100101101101011101100011"), -- 0.0184133 + 6.50314e-39 = 0.0184133
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010101110010101111101", b"10000000000010101110010101111101"), -- 0 + -1.00068e-39 = -1.00068e-39
	(b"01101001010011000010010000100001", b"00000000000000000000000000000000"),
	(b"10000000000010011101010110101111", b"01101001010011000010010000100001"), -- 1.54245e+25 + -9.03175e-40 = 1.54245e+25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111010001111001000110", b"11111111100000000000000000000000"), -- -inf + 5.61283e-39 = -inf
	(b"11101001001000010000100101000010", b"00000000000000000000000000000000"),
	(b"10000000010010111111010101111001", b"11101001001000010000100101000010"), -- -1.21675e+25 + -6.97572e-39 = -1.21675e+25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011010101001111110100000", b"11111111100000000000000000000000"), -- -inf + 9.79183e-39 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011100111010101011101011", b"00000000011100111010101011101011"), -- 0 + 1.06224e-38 = 1.06224e-38
	(b"10000000000000000000000001110011", b"00000000000000000000000000000000"),
	(b"00000000010010000100001010111101", b"00000000010010000100001001001010"), -- -1.61149e-43 + 6.6361e-39 = 6.63594e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001011011100110010101110", b"11111111100000000000000000000000"), -- -inf + -4.20602e-39 = -inf
	(b"00111110101001000000001000001001", b"00000000000000000000000000000000"),
	(b"10000000011010000100001110001001", b"00111110101001000000001000001001"), -- 0.320328 + -9.57512e-39 = 0.320328
	(b"00000000000000000000100010111000", b"00000000000000000000000000000000"),
	(b"00000000011000001110101101101111", b"00000000011000001111010000100111"), -- 3.1277e-42 + 8.90067e-39 = 8.90379e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001011100010101010010", b"00000000010001011100010101010010"), -- -0 + 6.40743e-39 = 6.40743e-39
	(b"10011010010010111100010101011011", b"00000000000000000000000000000000"),
	(b"00000000010111111001011010010100", b"10011010010010111100010101011011"), -- -4.21388e-23 + 8.77839e-39 = -4.21388e-23
	(b"10000000000000000011110100101001", b"00000000000000000000000000000000"),
	(b"00000000001111101011010100110111", b"00000000001111100111100000001110"), -- -2.19401e-41 + 5.75881e-39 = 5.73687e-39
	(b"10100100111100011010110011001111", b"00000000000000000000000000000000"),
	(b"00000000000110010000110000010001", b"10100100111100011010110011001111"), -- -1.0481e-16 + 2.30022e-39 = -1.0481e-16
	(b"01100111011101011111111000101101", b"00000000000000000000000000000000"),
	(b"00000000011101010101101000010000", b"01100111011101011111111000101101"), -- 1.16167e+24 + 1.07771e-38 = 1.16167e+24
	(b"00110111101101100111111010100001", b"00000000000000000000000000000000"),
	(b"00000000011010110100110010100010", b"00110111101101100111111010100001"), -- 2.17551e-05 + 9.85389e-39 = 2.17551e-05
	(b"00100111010100110000100101011111", b"00000000000000000000000000000000"),
	(b"10000000010100011111111010111000", b"00100111010100110000100101011111"), -- 2.92872e-15 + -7.53005e-39 = 2.92872e-15
	(b"00000000000000000010001001001000", b"00000000000000000000000000000000"),
	(b"10000000000101111101100010011001", b"10000000000101111011011001010001"), -- 1.22978e-41 + -2.18992e-39 = -2.17762e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101100010010000000000", b"00000000011101100010010000000000"), -- -0 + 1.08495e-38 = 1.08495e-38
	(b"01110100110000010110011100010001", b"00000000000000000000000000000000"),
	(b"00000000001011101101010000010011", b"01110100110000010110011100010001"), -- 1.22583e+32 + 4.30051e-39 = 1.22583e+32
	(b"00000000000000000000000000000010", b"00000000000000000000000000000000"),
	(b"00000000011101111100000110011001", b"00000000011101111100000110011011"), -- 2.8026e-45 + 1.09979e-38 = 1.09979e-38
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111001001100111000110", b"01111111100000000000000000000000"), -- inf + 5.56529e-39 = inf
	(b"10000000000010100100110011110010", b"00000000000000000000000000000000"),
	(b"00000000001001010100100011001000", b"00000000000110101111101111010110"), -- -9.45958e-40 + 3.42402e-39 = 2.47806e-39
	(b"10000000000000101000110000010100", b"00000000000000000000000000000000"),
	(b"00000000001000110000010110110011", b"00000000001000000111100110011111"), -- -2.33922e-40 + 3.21629e-39 = 2.98237e-39
	(b"11011101010111011001100001111011", b"00000000000000000000000000000000"),
	(b"00000000001010100001011000000110", b"11011101010111011001100001111011"), -- -9.97978e+17 + 3.86499e-39 = -9.97978e+17
	(b"10000111001000010000100111110011", b"00000000000000000000000000000000"),
	(b"00000000011000111100010100010011", b"10000111001000010000011011010101"), -- -1.21152e-34 + 9.16241e-39 = -1.21143e-34
	(b"11010100011000000100100010111000", b"00000000000000000000000000000000"),
	(b"00000000001001110101100001011111", b"11010100011000000100100010111000"), -- -3.85317e+12 + 3.61329e-39 = -3.85317e+12
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010100000001010101101011", b"10000000010100000001010101101011"), -- 0 + -7.35452e-39 = -7.35452e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011011001010001100000111", b"10000000011011001010001100000111"), -- 0 + -9.97672e-39 = -9.97672e-39
	(b"10000000000000000000000000001101", b"00000000000000000000000000000000"),
	(b"00000000000000010000100000110001", b"00000000000000010000100000100100"), -- -1.82169e-44 + 9.4774e-41 = 9.47558e-41
	(b"11111101000010001111010001011111", b"00000000000000000000000000000000"),
	(b"00000000000110110011001100000111", b"11111101000010001111010001011111"), -- -1.13777e+37 + 2.49786e-39 = -1.13777e+37
	(b"00011110011001110110010011010011", b"00000000000000000000000000000000"),
	(b"10000000000001011100001110111100", b"00011110011001110110010011010011"), -- 1.22499e-20 + -5.29394e-40 = 1.22499e-20
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"10000000000001101011110011110011", b"10000000000001101011110011110100"), -- -1.4013e-45 + -6.18795e-40 = -6.18797e-40
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110001110111100010000", b"00000000000110001110111100010000"), -- -0 + 2.28981e-39 = 2.28981e-39
	(b"01010110000001111111010110101101", b"00000000000000000000000000000000"),
	(b"00000000011111010110101101001011", b"01010110000001111111010110101101"), -- 3.73723e+13 + 1.15179e-38 = 3.73723e+13
	(b"00101010100000010100001010111100", b"00000000000000000000000000000000"),
	(b"00000000001111101100011111101111", b"00101010100000010100001010111100"), -- 2.29613e-13 + 5.76552e-39 = 2.29613e-13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000001011001101101000", b"01111111100000000000000000000000"), -- inf + 6.43588e-41 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111110110110101110100", b"10000000010111110110110101110100"), -- -0 + -8.76364e-39 = -8.76364e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001111010010100100101001", b"10000000001111010010100100101001"), -- -0 + -5.61673e-39 = -5.61673e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010001001110101010010100", b"01111111100000000000000000000000"), -- inf + -6.32896e-39 = inf
	(b"00000000000000000000000001011011", b"00000000000000000000000000000000"),
	(b"00000000000101010111000010000010", b"00000000000101010111000011011101"), -- 1.27518e-43 + 1.96891e-39 = 1.96903e-39
	(b"11110110000100111110101110010001", b"00000000000000000000000000000000"),
	(b"10000000010101000001111010011000", b"11110110000100111110101110010001"), -- -7.50044e+32 + -7.72516e-39 = -7.50044e+32
	(b"11101000100000011111010011010011", b"00000000000000000000000000000000"),
	(b"00000000000010010001010110110011", b"11101000100000011111010011010011"), -- -4.90961e+24 + 8.34304e-40 = -4.90961e+24
	(b"00011101001101011010111010001101", b"00000000000000000000000000000000"),
	(b"00000000001010011101000101110001", b"00011101001101011010111010001101"), -- 2.40454e-21 + 3.84039e-39 = 2.40454e-21
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010010100001011100101", b"11111111100000000000000000000000"), -- -inf + 8.50517e-40 = -inf
	(b"00000000000000000010100101000011", b"00000000000000000000000000000000"),
	(b"10000000011100110101001101010011", b"10000000011100110010101000010000"), -- 1.48019e-41 + -1.0591e-38 = -1.05762e-38
	(b"11100001100100110000011000001111", b"00000000000000000000000000000000"),
	(b"00000000010000111011001110000011", b"11100001100100110000011000001111"), -- -3.39013e+20 + 6.21737e-39 = -3.39013e+20
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001010001110011111110", b"01111111100000000000000000000000"), -- inf + -9.28579e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010111010000011111001", b"11111111100000000000000000000000"), -- -inf + 4.00667e-39 = -inf
	(b"10000000000010001011110100101101", b"00000000000000000000000000000000"),
	(b"00000000000011001011111010100000", b"00000000000001000000000101110011"), -- -8.02547e-40 + 1.17041e-39 = 3.67862e-40
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010011000001001101111", b"10000000000010011000001001101111"), -- 0 + -8.7331e-40 = -8.7331e-40
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010101100101110001100001", b"10000000010101100101110001100001"), -- 0 + -7.93099e-39 = -7.93099e-39
	(b"11110111101011111000000111100111", b"00000000000000000000000000000000"),
	(b"00000000001000111000101110011110", b"11110111101011111000000111100111"), -- -7.11943e+33 + 3.26433e-39 = -7.11943e+33
	(b"00001101100001101010111110100011", b"00000000000000000000000000000000"),
	(b"10000000011101111111101010011110", b"00001101100001101010111110100011"), -- 8.30067e-31 + -1.10183e-38 = 8.30067e-31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111010011110110010111", b"11111111100000000000000000000000"), -- -inf + -8.5628e-39 = -inf
	(b"00011010111100001111001001001001", b"00000000000000000000000000000000"),
	(b"10000000001001000100100111011110", b"00011010111100001111001001001001"), -- 9.96531e-23 + -3.33258e-39 = 9.96531e-23
	(b"10101101101111111010110001100110", b"00000000000000000000000000000000"),
	(b"10000000000110010111101001100110", b"10101101101111111010110001100110"), -- -2.17907e-11 + -2.3398e-39 = -2.17907e-11
	(b"01000001010000001011110101110110", b"00000000000000000000000000000000"),
	(b"00000000010010000101010110011001", b"01000001010000001011110101110110"), -- 12.0463 + 6.64286e-39 = 12.0463
	(b"11111100111100010000001001101110", b"00000000000000000000000000000000"),
	(b"00000000011110101001100111101010", b"11111100111100010000001001101110"), -- -1.00111e+37 + 1.12591e-38 = -1.00111e+37
	(b"01110101001011000000001111111110", b"00000000000000000000000000000000"),
	(b"10000000011001011110011000010110", b"01110101001011000000001111111110"), -- 2.18056e+32 + -9.35792e-39 = 2.18056e+32
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110111010010111111010", b"11111111100000000000000000000000"), -- -inf + -8.41657e-39 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010100101100011011010110", b"00000000010100101100011011010110"), -- -0 + 7.60184e-39 = 7.60184e-39
	(b"01110010010101010111110011111111", b"00000000000000000000000000000000"),
	(b"10000000010000100101101100110101", b"01110010010101010111110011111111"), -- 4.22857e+30 + -6.09386e-39 = 4.22857e+30
	(b"11011001101011100110001110100101", b"00000000000000000000000000000000"),
	(b"10000000011111010010101010001010", b"11011001101011100110001110100101"), -- -6.13578e+15 + -1.14947e-38 = -6.13578e+15
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011010100010010110110", b"00000000001011010100010010110110"), -- 0 + 4.15725e-39 = 4.15725e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001100000011101111011100", b"10000000001100000011101111011100"), -- -0 + -4.42958e-39 = -4.42958e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001111011101110100110111", b"10000000001111011101110100110111"), -- -0 + -5.68132e-39 = -5.68132e-39
	(b"00101101111100110100010111101101", b"00000000000000000000000000000000"),
	(b"00000000010011010110001100101000", b"00101101111100110100010111101101"), -- 2.7657e-11 + 7.1069e-39 = 2.7657e-11
	(b"00101011100111000111101111010111", b"00000000000000000000000000000000"),
	(b"10000000011001111100110101111010", b"00101011100111000111101111010111"), -- 1.11188e-12 + -9.53277e-39 = 1.11188e-12
	(b"01010101100011111101010101010101", b"00000000000000000000000000000000"),
	(b"10000000000100100100000010111010", b"01010101100011111101010101010101"), -- 1.97683e+13 + -1.67626e-39 = 1.97683e+13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010011111111011111101100", b"01111111100000000000000000000000"), -- inf + 7.34394e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000011000110101001010", b"01111111100000000000000000000000"), -- inf + -8.95873e-39 = inf
	(b"11111101111010101000110110000000", b"00000000000000000000000000000000"),
	(b"10000000010000111001010101010101", b"11111101111010101000110110000000"), -- -3.89718e+37 + -6.20655e-39 = -3.89718e+37
	(b"00101100101111110100110011001011", b"00000000000000000000000000000000"),
	(b"10000000000100111000100101010001", b"00101100101111110100110011001011"), -- 5.43707e-12 + -1.79413e-39 = 5.43707e-12
	(b"01110110000001100111110001011000", b"00000000000000000000000000000000"),
	(b"00000000000000111110100001111101", b"01110110000001100111110001011000"), -- 6.81924e+32 + 3.58908e-40 = 6.81924e+32
	(b"10111001110001001000111000010000", b"00000000000000000000000000000000"),
	(b"10000000000101001101000010001010", b"10111001110001001000111000010000"), -- -0.000374899 + -1.91152e-39 = -0.000374899
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001111001110111010101", b"11111111100000000000000000000000"), -- -inf + 6.57694e-39 = -inf
	(b"00110001101010110001001100101111", b"00000000000000000000000000000000"),
	(b"00000000011101111001100011000010", b"00110001101010110001001100101111"), -- 4.97894e-09 + 1.09832e-38 = 4.97894e-09
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000101011111010011111", b"11111111100000000000000000000000"), -- -inf + 2.52053e-40 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010000000001110111100100", b"01111111100000000000000000000000"), -- inf + -5.88819e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011000000101110101101101", b"00000000011000000101110101101101"), -- 0 + 8.84972e-39 = 8.84972e-39
	(b"00111111010111111110010000100110", b"00000000000000000000000000000000"),
	(b"00000000000101000011111111011111", b"00111111010111111110010000100110"), -- 0.874575 + 1.85962e-39 = 0.874575
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001111111010011011000", b"11111111100000000000000000000000"), -- -inf + 6.60815e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010110001110010110001", b"01111111100000000000000000000000"), -- inf + 1.02048e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101000101111000011111", b"11111111100000000000000000000000"), -- -inf + 1.06867e-38 = -inf
	(b"00001001010110010011100110011000", b"00000000000000000000000000000000"),
	(b"10000000011011111100010101100110", b"00001001010110010011100101100000"), -- 2.61475e-33 + -1.02646e-38 = 2.61474e-33
	(b"10000000000101001101100010110011", b"00000000000000000000000000000000"),
	(b"00000000011011000011111100100101", b"00000000010101110110011001110010"), -- -1.91445e-39 + 9.94089e-39 = 8.02644e-39
	(b"01111111000111110100100001110101", b"00000000000000000000000000000000"),
	(b"10000000010100000010100011110110", b"01111111000111110100100001110101"), -- 2.11723e+38 + -7.36153e-39 = 2.11723e+38
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011111101001011001110", b"11111111100000000000000000000000"), -- -inf + 1.45315e-39 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101110110011011110111", b"10000000001101110110011011110111"), -- -0 + -5.08789e-39 = -5.08789e-39
	(b"00100101000100001000000100100100", b"00000000000000000000000000000000"),
	(b"00000000000110011111110101101010", b"00100101000100001000000100100100"), -- 1.25338e-16 + 2.3868e-39 = 1.25338e-16
	(b"10100010001000101011111001000010", b"00000000000000000000000000000000"),
	(b"10000000011111010111111110011001", b"10100010001000101011111001000010"), -- -2.20558e-18 + -1.15252e-38 = -2.20558e-18
	(b"11011011001101001000110101001010", b"00000000000000000000000000000000"),
	(b"10000000001001000000000000111000", b"11011011001101001000110101001010"), -- -5.08208e+16 + -3.30616e-39 = -5.08208e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011001111010111010011", b"11111111100000000000000000000000"), -- -inf + 1.00064e-38 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011100100100100111101010", b"00000000011100100100100111101010"), -- 0 + 1.04958e-38 = 1.04958e-38
	(b"00000110100011001101001100010110", b"00000000000000000000000000000000"),
	(b"10000000010110011100001100100000", b"00000110100011001100110101111010"), -- 5.29723e-35 + -8.24336e-39 = 5.29641e-35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000110010000000100101000", b"11111111100000000000000000000000"), -- -inf + -2.2963e-39 = -inf
	(b"10010100111000010110010000110010", b"00000000000000000000000000000000"),
	(b"10000000001110010010000110100110", b"10010100111000010110010000110010"), -- -2.27587e-26 + -5.24669e-39 = -2.27587e-26
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001000011000010111011", b"01111111100000000000000000000000"), -- inf + -3.32356e-39 = inf
	(b"00100011000110100110000100100010", b"00000000000000000000000000000000"),
	(b"10000000011110111110011100100111", b"00100011000110100110000100100010"), -- 8.36893e-18 + -1.13787e-38 = 8.36893e-18
	(b"00000000000000000110110111010111", b"00000000000000000000000000000000"),
	(b"10000000000111000101000001011010", b"10000000000110111110001010000011"), -- 3.94031e-41 + -2.60022e-39 = -2.56082e-39
	(b"00101110001110001101010011111011", b"00000000000000000000000000000000"),
	(b"00000000011100100000100001011110", b"00101110001110001101010011111011"), -- 4.20259e-11 + 1.04722e-38 = 4.20259e-11
	(b"11011111101000011000011111101000", b"00000000000000000000000000000000"),
	(b"10000000000110101010011000000110", b"11011111101000011000011111101000"), -- -2.32791e+19 + -2.44728e-39 = -2.32791e+19
	(b"11011010111111111101100100011101", b"00000000000000000000000000000000"),
	(b"10000000001011101110000001011011", b"11011010111111111101100100011101"), -- -3.60074e+16 + -4.30492e-39 = -3.60074e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011001101111101110110", b"11111111100000000000000000000000"), -- -inf + -1.18219e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001100011110011110101", b"11111111100000000000000000000000"), -- -inf + 6.45035e-39 = -inf
	(b"10000000000000000000000000000101", b"00000000000000000000000000000000"),
	(b"00000000011001010010010110110101", b"00000000011001010010010110110000"), -- -7.00649e-45 + 9.28891e-39 = 9.2889e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001010101000101100110", b"01111111100000000000000000000000"), -- inf + 9.30459e-39 = inf
	(b"00001011010111000111101100110101", b"00000000000000000000000000000000"),
	(b"10000000001101101111100011001011", b"00001011010111000111101100110011"), -- 4.24631e-32 + -5.04837e-39 = 4.24631e-32
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011001100101110000101", b"00000000001011001100101110000101"), -- 0 + 4.11377e-39 = 4.11377e-39
	(b"00111110101001101010101111010000", b"00000000000000000000000000000000"),
	(b"00000000001111100100011101010111", b"00111110101001101010101111010000"), -- 0.32553 + 5.71939e-39 = 0.32553
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011100010100101010100", b"01111111100000000000000000000000"), -- inf + 1.01167e-38 = inf
	(b"10011000011011010111010011000110", b"00000000000000000000000000000000"),
	(b"00000000011100111000100011111000", b"10011000011011010111010011000110"), -- -3.06905e-24 + 1.06102e-38 = -3.06905e-24
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000011010100000011", b"00000000000000000011010100000011"), -- 0 + 1.9017e-41 = 1.9017e-41
	(b"01000011011111111001111100100011", b"00000000000000000000000000000000"),
	(b"00000000001110011011101011011000", b"01000011011111111001111100100011"), -- 255.622 + 5.30165e-39 = 255.622
	(b"11001111100111100101010101100000", b"00000000000000000000000000000000"),
	(b"10000000000110110000011110100000", b"11001111100111100101010101100000"), -- -5.31279e+09 + -2.48229e-39 = -5.31279e+09
	(b"01111011100000110100011111111000", b"00000000000000000000000000000000"),
	(b"00000000010010001111011110100000", b"01111011100000110100011111111000"), -- 1.3633e+36 + 6.70099e-39 = 1.3633e+36
	(b"10001000101100010010110100101101", b"00000000000000000000000000000000"),
	(b"10000000011000111100100001110111", b"10001000101100010010110110010001"), -- -1.06634e-33 + -9.16363e-39 = -1.06635e-33
	(b"00101001000110101011010000010000", b"00000000000000000000000000000000"),
	(b"00000000001101111101110011000110", b"00101001000110101011010000010000"), -- 3.4351e-14 + 5.13015e-39 = 3.4351e-14
	(b"01101010101001001110101110011101", b"00000000000000000000000000000000"),
	(b"10000000000001101110101111000001", b"01101010101001001110101110011101"), -- 9.96882e+25 + -6.35586e-40 = 9.96882e+25
	(b"11010011000001000000111111110110", b"00000000000000000000000000000000"),
	(b"00000000001001110010000001010001", b"11010011000001000000111111110110"), -- -5.67203e+11 + 3.59318e-39 = -5.67203e+11
	(b"00101101101011110101111010011001", b"00000000000000000000000000000000"),
	(b"00000000010011100000100001011010", b"00101101101011110101111010011001"), -- 1.99372e-11 + 7.16616e-39 = 1.99372e-11
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001100111010100011101", b"11111111100000000000000000000000"), -- -inf + -9.40923e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110101111011000001110", b"11111111100000000000000000000000"), -- -inf + 2.47599e-39 = -inf
	(b"10010011010001110111001110111011", b"00000000000000000000000000000000"),
	(b"10000000000010000111001100110011", b"10010011010001110111001110111011"), -- -2.51744e-27 + -7.7601e-40 = -2.51744e-27
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000010111011100000001111", b"01111111100000000000000000000000"), -- inf + 1.07622e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110111101100111010101", b"01111111100000000000000000000000"), -- inf + 5.49644e-39 = inf
	(b"00010101111100001010110000100110", b"00000000000000000000000000000000"),
	(b"10000000010110011001101010011000", b"00010101111100001010110000100110"), -- 9.72068e-26 + -8.22882e-39 = 9.72068e-26
	(b"01110110110000010010111011101001", b"00000000000000000000000000000000"),
	(b"10000000011110011000111110011111", b"01110110110000010010111011101001"), -- 1.95911e+33 + -1.11636e-38 = 1.95911e+33
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000111100001000010110100", b"10000000000111100001000010110100"), -- -0 + -2.76106e-39 = -2.76106e-39
	(b"01101011101001010110101001101111", b"00000000000000000000000000000000"),
	(b"10000000010101010000100000010000", b"01101011101001010110101001101111"), -- 3.99951e+26 + -7.80891e-39 = 3.99951e+26
	(b"11100000001110001111001000100110", b"00000000000000000000000000000000"),
	(b"00000000010101010110011110001101", b"11100000001110001111001000100110"), -- -5.3307e+19 + 7.84316e-39 = -5.3307e+19
	(b"11100011000000010111001110100101", b"00000000000000000000000000000000"),
	(b"10000000010000000010010111100111", b"11100011000000010111001110100101"), -- -2.38796e+21 + -5.89107e-39 = -2.38796e+21
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001110111010100010101", b"01111111100000000000000000000000"), -- inf + 6.56232e-39 = inf
	(b"00001110111000111011000000011100", b"00000000000000000000000000000000"),
	(b"00000000001000011001100010101001", b"00001110111000111011000000011100"), -- 5.61294e-30 + 3.08534e-39 = 5.61294e-30
	(b"11101011011001110011110111010010", b"00000000000000000000000000000000"),
	(b"00000000000111001110101000110010", b"11101011011001110011110111010010"), -- -2.79554e+26 + 2.65541e-39 = -2.79554e+26
	(b"11110001110111001011011111001011", b"00000000000000000000000000000000"),
	(b"10000000001110101001111100110001", b"11110001110111001011011111001011"), -- -2.18588e+30 + -5.38357e-39 = -2.18588e+30
	(b"10011011100001101100001110010010", b"00000000000000000000000000000000"),
	(b"00000000001011001111100011111101", b"10011011100001101100001110010010"), -- -2.22948e-22 + 4.13008e-39 = -2.22948e-22
	(b"00010011110000111011010010111100", b"00000000000000000000000000000000"),
	(b"00000000010111010011000001001110", b"00010011110000111011010010111100"), -- 4.94031e-27 + 8.55803e-39 = 4.94031e-27
	(b"00101111001100010100011110011001", b"00000000000000000000000000000000"),
	(b"10000000000011000101011101011111", b"00101111001100010100011110011001"), -- 1.61235e-10 + -1.13337e-39 = 1.61235e-10
	(b"10000000000000000000000011110001", b"00000000000000000000000000000000"),
	(b"10000000001111001001000011101100", b"10000000001111001001000111011101"), -- -3.37713e-43 + -5.56212e-39 = -5.56246e-39
	(b"00100100100010101100011011000111", b"00000000000000000000000000000000"),
	(b"10000000010011010001010100011011", b"00100100100010101100011011000111"), -- 6.01847e-17 + -7.0789e-39 = 6.01847e-17
	(b"10010110011010111111001110001101", b"00000000000000000000000000000000"),
	(b"10000000011100111000111010000011", b"10010110011010111111001110001101"), -- -1.906e-25 + -1.06122e-38 = -1.906e-25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011011100001000101001", b"11111111100000000000000000000000"), -- -inf + 1.26351e-39 = -inf
	(b"11000011010000001110010100010011", b"00000000000000000000000000000000"),
	(b"10000000010110110101101000011101", b"11000011010000001110010100010011"), -- -192.895 + -8.38936e-39 = -192.895
	(b"11111100010010010110110111111101", b"00000000000000000000000000000000"),
	(b"00000000010101001101100110000001", b"11111100010010010110110111111101"), -- -4.18353e+36 + 7.79221e-39 = -4.18353e+36
	(b"00000000000000000010100111000000", b"00000000000000000000000000000000"),
	(b"10000000011111110010101101101111", b"10000000011111110000000110101111"), -- 1.49771e-41 + -1.16787e-38 = -1.16637e-38
	(b"00000000000000000000000000100100", b"00000000000000000000000000000000"),
	(b"00000000010001100000011000011110", b"00000000010001100000011001000010"), -- 5.04467e-44 + 6.43068e-39 = 6.43073e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001110110000111010111", b"11111111100000000000000000000000"), -- -inf + 6.77947e-40 = -inf
	(b"00101000011100110010101011000010", b"00000000000000000000000000000000"),
	(b"10000000011000111100010111000100", b"00101000011100110010101011000010"), -- 1.34985e-14 + -9.16266e-39 = 1.34985e-14
	(b"01010011010000011000101010000010", b"00000000000000000000000000000000"),
	(b"10000000011010011001110100100010", b"01010011010000011000101010000010"), -- 8.31252e+11 + -9.6991e-39 = 8.31252e+11
	(b"10111111011000101110100110101010", b"00000000000000000000000000000000"),
	(b"00000000000100001110101001110110", b"10111111011000101110100110101010"), -- -0.886378 + 1.55348e-39 = -0.886378
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001001000101110010101101", b"01111111100000000000000000000000"), -- inf + 3.33932e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011000101010110001100", b"00000000001011000101010110001100"), -- 0 + 4.07145e-39 = 4.07145e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101101000100011010100", b"10000000011101101000100011010100"), -- -0 + -1.08857e-38 = -1.08857e-38
	(b"11010111011110101111001101101100", b"00000000000000000000000000000000"),
	(b"00000000000111011111101110000111", b"11010111011110101111001101101100"), -- -2.75923e+14 + 2.75346e-39 = -2.75923e+14
	(b"10111101100001010010001100010110", b"00000000000000000000000000000000"),
	(b"10000000000101100000101001111111", b"10111101100001010010001100010110"), -- -0.0650083 + -2.02415e-39 = -0.0650083
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110110110010001110000", b"11111111100000000000000000000000"), -- -inf + 2.51559e-39 = -inf
	(b"10001000011110101111010100101110", b"00000000000000000000000000000000"),
	(b"00000000001011110100011111100000", b"10001000011110101111010011001111"), -- -7.55198e-34 + 4.34205e-39 = -7.55194e-34
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000101011110010010001001", b"01111111100000000000000000000000"), -- inf + 2.01053e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010010011011010100100", b"11111111100000000000000000000000"), -- -inf + 3.78486e-39 = -inf
	(b"11100110011010000001110011010111", b"00000000000000000000000000000000"),
	(b"00000000010111001011110101111110", b"11100110011010000001110011010111"), -- -2.7403e+23 + 8.51684e-39 = -2.7403e+23
	(b"00010101110011001010101010010100", b"00000000000000000000000000000000"),
	(b"00000000000011000111011000000100", b"00010101110011001010101010010100"), -- 8.26641e-26 + 1.14436e-39 = 8.26641e-26
	(b"11010001001011110100010101010100", b"00000000000000000000000000000000"),
	(b"10000000011010101110111010100011", b"11010001001011110100010101010100"), -- -4.70489e+10 + -9.82017e-39 = -4.70489e+10
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010111111101001001100", b"10000000000010111111101001001100"), -- -0 + -1.09998e-39 = -1.09998e-39
	(b"11110100011001001011101111111100", b"00000000000000000000000000000000"),
	(b"00000000010001001110011110000011", b"11110100011001001011101111111100"), -- -7.24888e+31 + 6.32786e-39 = -7.24888e+31
	(b"00001111111001011011000010110100", b"00000000000000000000000000000000"),
	(b"00000000000101111100101101111010", b"00001111111001011011000010110100"), -- 2.26492e-29 + 2.18521e-39 = 2.26492e-29
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101101100110100101001", b"00000000011101101100110100101001"), -- 0 + 1.09102e-38 = 1.09102e-38
	(b"01001101100100001010100111111000", b"00000000000000000000000000000000"),
	(b"00000000011011010100110111100101", b"01001101100100001010100111111000"), -- 3.03382e+08 + 1.0038e-38 = 3.03382e+08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010111010111111000000110", b"01111111100000000000000000000000"), -- inf + 8.58591e-39 = inf
	(b"10011000001011010110110010111000", b"00000000000000000000000000000000"),
	(b"10000000000010010011001101110010", b"10011000001011010110110010111000"), -- -2.24146e-24 + -8.44975e-40 = -2.24146e-24
	(b"01001010010001101111110111110001", b"00000000000000000000000000000000"),
	(b"10000000010000110010011010010000", b"01001010010001101111110111110001"), -- 3.26028e+06 + -6.16681e-39 = 3.26028e+06
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111111111000001111110", b"11111111100000000000000000000000"), -- -inf + -8.81064e-39 = -inf
	(b"11100110010100110111011101111111", b"00000000000000000000000000000000"),
	(b"00000000010011010011000101111110", b"11100110010100110111011101111111"), -- -2.49656e+23 + 7.08909e-39 = -2.49656e+23
	(b"11101100101011011111101010100111", b"00000000000000000000000000000000"),
	(b"00000000000100011001110010010111", b"11101100101011011111101010100111"), -- -1.68262e+27 + 1.61738e-39 = -1.68262e+27
	(b"11110000010111011101001000111101", b"00000000000000000000000000000000"),
	(b"10000000000110010100010001101011", b"11110000010111011101001000111101"), -- -2.74601e+29 + -2.32043e-39 = -2.74601e+29
	(b"00000111101001011010111011110111", b"00000000000000000000000000000000"),
	(b"00000000011101110011101010110101", b"00000111101001011011000011010100"), -- 2.49293e-34 + 1.09495e-38 = 2.49304e-34
	(b"00111110010111011111110101111101", b"00000000000000000000000000000000"),
	(b"10000000011111001000100010000100", b"00111110010111011111110101111101"), -- 0.216787 + -1.14366e-38 = 0.216787
	(b"00101101100001100001010110010010", b"00000000000000000000000000000000"),
	(b"10000000001111101110001001100001", b"00101101100001100001010110010010"), -- 1.52436e-11 + -5.77501e-39 = 1.52436e-11
	(b"00000010111011101100111110001000", b"00000000000000000000000000000000"),
	(b"00000000000101110011010010101111", b"00000010111100000100001011010011"), -- 3.50901e-37 + 2.13112e-39 = 3.53032e-37
	(b"00111000010000011010100101000110", b"00000000000000000000000000000000"),
	(b"00000000001001010111111110111110", b"00111000010000011010100101000110"), -- 4.61724e-05 + 3.44374e-39 = 4.61724e-05
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110111001000010110000", b"00000000000110111001000010110000"), -- 0 + 2.53146e-39 = 2.53146e-39
	(b"01010101001110010111001011001000", b"00000000000000000000000000000000"),
	(b"00000000011100001111010110010111", b"01010101001110010111001011001000"), -- 1.27439e+13 + 1.03737e-38 = 1.27439e+13
	(b"01101001110000100011110011111111", b"00000000000000000000000000000000"),
	(b"00000000011000010110001010000001", b"01101001110000100011110011111111"), -- 2.93525e+25 + 8.94338e-39 = 2.93525e+25
	(b"11001110101101000100001100011000", b"00000000000000000000000000000000"),
	(b"10000000000101010101000001111000", b"11001110101101000100001100011000"), -- -1.51215e+09 + -1.95741e-39 = -1.51215e+09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001000001111100111010", b"01111111100000000000000000000000"), -- inf + -9.19475e-39 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011110111110001011111010", b"00000000011110111110001011111010"), -- -0 + 1.13772e-38 = 1.13772e-38
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110110011101011000101", b"11111111100000000000000000000000"), -- -inf + 5.43938e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001100101000100110110001", b"11111111100000000000000000000000"), -- -inf + -4.64117e-39 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110010010010110101100", b"00000000010110010010010110101100"), -- 0 + 8.18687e-39 = 8.18687e-39
	(b"00101001001000000101101111000011", b"00000000000000000000000000000000"),
	(b"00000000000000110000000110110110", b"00101001001000000101101111000011"), -- 3.56067e-14 + 2.7612e-40 = 3.56067e-14
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001000110011111110000", b"11111111100000000000000000000000"), -- -inf + -3.34336e-39 = -inf
	(b"10111111100001110111110000101101", b"00000000000000000000000000000000"),
	(b"10000000001100010100001110011100", b"10111111100001110111110000101101"), -- -1.05848 + -4.52419e-39 = -1.05848
	(b"10011011111000011011110001111001", b"00000000000000000000000000000000"),
	(b"00000000011100001111011101001100", b"10011011111000011011110001111001"), -- -3.73449e-22 + 1.03743e-38 = -3.73449e-22
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110010111011001011000", b"01111111100000000000000000000000"), -- inf + 5.27708e-39 = inf
	(b"10011011111010001100010011111111", b"00000000000000000000000000000000"),
	(b"00000000011110010110101100000000", b"10011011111010001100010011111111"), -- -3.85085e-22 + 1.11505e-38 = -3.85085e-22
	(b"01010001111110000011010000101111", b"00000000000000000000000000000000"),
	(b"10000000000000100001101010101001", b"01010001111110000011010000101111"), -- 1.33253e+11 + -1.93235e-40 = 1.33253e+11
	(b"10111110000101100111100111101110", b"00000000000000000000000000000000"),
	(b"00000000000100110001000111110011", b"10111110000101100111100111101110"), -- -0.146949 + 1.75131e-39 = -0.146949
	(b"00111110100000001000010000100011", b"00000000000000000000000000000000"),
	(b"10000000010000111110111001000010", b"00111110100000001000010000100011"), -- 0.251008 + -6.23845e-39 = 0.251008
	(b"00100111100010100001010111101100", b"00000000000000000000000000000000"),
	(b"10000000010010011001010101110010", b"00100111100010100001010111101100"), -- 3.83265e-15 + -6.7576e-39 = 3.83265e-15
	(b"11101111110100101010110100001111", b"00000000000000000000000000000000"),
	(b"10000000011101110001100111101000", b"11101111110100101010110100001111"), -- -1.30402e+29 + -1.09377e-38 = -1.30402e+29
	(b"00111111010110101000100011001000", b"00000000000000000000000000000000"),
	(b"10000000011110100000010111011001", b"00111111010110101000100011001000"), -- 0.85365 + -1.1206e-38 = 0.85365
	(b"00001101010100010100010010001001", b"00000000000000000000000000000000"),
	(b"10000000001000100100010101101110", b"00001101010100010100010010001001"), -- 6.44856e-31 + -3.14731e-39 = 6.44856e-31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010101100010101101100", b"00000000001010101100010101101100"), -- -0 + 3.92791e-39 = 3.92791e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111111101011010000110", b"01111111100000000000000000000000"), -- inf + 5.86259e-39 = inf
	(b"00101101100001001101110001001010", b"00000000000000000000000000000000"),
	(b"10000000010110010110001000011001", b"00101101100001001101110001001010"), -- 1.51045e-11 + -8.20855e-39 = 1.51045e-11
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110101000111011010100", b"10000000001110101000111011010100"), -- -0 + -5.3777e-39 = -5.3777e-39
	(b"11001110100100110000100011100100", b"00000000000000000000000000000000"),
	(b"00000000010011011110001101111001", b"11001110100100110000100011100100"), -- -1.23342e+09 + 7.15294e-39 = -1.23342e+09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011000000001110111011101", b"01111111100000000000000000000000"), -- inf + 8.82692e-39 = inf
	(b"11100000101011011101100110110011", b"00000000000000000000000000000000"),
	(b"00000000011000101101001100110000", b"11100000101011011101100110110011"), -- -1.00218e+20 + 9.07564e-39 = -1.00218e+20
	(b"11000100010100010110001001101011", b"00000000000000000000000000000000"),
	(b"10000000010000101111110011001001", b"11000100010100010110001001101011"), -- -837.538 + -6.15182e-39 = -837.538
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000000111000100110011", b"10000000011000000111000100110011"), -- 0 + -8.85682e-39 = -8.85682e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111111001101000010110", b"01111111100000000000000000000000"), -- inf + 2.90218e-39 = inf
	(b"00101011001011111001010001111000", b"00000000000000000000000000000000"),
	(b"10000000000010011111100101011101", b"00101011001011111001010001111000"), -- 6.23785e-13 + -9.15974e-40 = 6.23785e-13
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100010001110010110101", b"10000000011100010001110010110101"), -- -0 + -1.03877e-38 = -1.03877e-38
	(b"11100000001010110010011111000100", b"00000000000000000000000000000000"),
	(b"10000000000110110100000011111010", b"11100000001010110010011111000100"), -- -4.93322e+19 + -2.50287e-39 = -4.93322e+19
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101000000100111110011", b"10000000001101000000100111110011"), -- -0 + -4.77901e-39 = -4.77901e-39
	(b"00000000000000000000000000000100", b"00000000000000000000000000000000"),
	(b"10000000011001010001101100111101", b"10000000011001010001101100111001"), -- 5.60519e-45 + -9.28516e-39 = -9.28515e-39
	(b"10010100100001011111000101001000", b"00000000000000000000000000000000"),
	(b"00000000001111100100000110101010", b"10010100100001011111000101001000"), -- -1.35247e-26 + 5.71736e-39 = -1.35247e-26
	(b"00101001100011100001010100011111", b"00000000000000000000000000000000"),
	(b"00000000010000011011011101101010", b"00101001100011100001010100011111"), -- 6.30973e-14 + 6.0351e-39 = 6.30973e-14
	(b"01111000100101111101010100111110", b"00000000000000000000000000000000"),
	(b"00000000000100111101001010110101", b"01111000100101111101010100111110"), -- 2.46363e+34 + 1.82046e-39 = 2.46363e+34
	(b"10010100100101101010101100101001", b"00000000000000000000000000000000"),
	(b"10000000010110111001101010101111", b"10010100100101101010101100101001"), -- -1.52136e-26 + -8.41252e-39 = -1.52136e-26
	(b"10011010110010101100011110010110", b"00000000000000000000000000000000"),
	(b"10000000000111101000000101111110", b"10011010110010101100011110010110"), -- -8.38677e-23 + -2.80152e-39 = -8.38677e-23
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010000011100001000010", b"01111111100000000000000000000000"), -- inf + 3.6936e-39 = inf
	(b"01011100100110001011111010010100", b"00000000000000000000000000000000"),
	(b"00000000010011100001111011011011", b"01011100100110001011111010010100"), -- 3.4395e+17 + 7.17424e-39 = 3.4395e+17
	(b"00001110101100101100110000101000", b"00000000000000000000000000000000"),
	(b"00000000011010000111101011001100", b"00001110101100101100110000101000"), -- 4.4077e-30 + 9.59494e-39 = 4.4077e-30
	(b"01100001010100111001110100001011", b"00000000000000000000000000000000"),
	(b"10000000010100101111111110111110", b"01100001010100111001110100001011"), -- 2.43974e+20 + -7.62225e-39 = 2.43974e+20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110110101010000100000", b"00000000001110110101010000100000"), -- -0 + 5.44847e-39 = 5.44847e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001010000110110101111", b"10000000001001010000110110101111"), -- -0 + -3.40282e-39 = -3.40282e-39
	(b"00001110011000000000100100000001", b"00000000000000000000000000000000"),
	(b"00000000000001001000011111100110", b"00001110011000000000100100000001"), -- 2.76145e-30 + 4.16093e-40 = 2.76145e-30
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010101110001010100011000", b"11111111100000000000000000000000"), -- -inf + -7.99726e-39 = -inf
	(b"11000001100011011000100001010000", b"00000000000000000000000000000000"),
	(b"00000000001000000100001001101110", b"11000001100011011000100001010000"), -- -17.6916 + 2.96257e-39 = -17.6916
	(b"00111101100110000000111101101011", b"00000000000000000000000000000000"),
	(b"10000000000011011101100001001101", b"00111101100110000000111101101011"), -- 0.0742482 + -1.27146e-39 = 0.0742482
	(b"10111010000000101000101000000001", b"00000000000000000000000000000000"),
	(b"00000000000010001011010111001101", b"10111010000000101000101000000001"), -- -0.000497967 + 7.99902e-40 = -0.000497967
	(b"10110000001101000100001010100000", b"00000000000000000000000000000000"),
	(b"10000000001110000000001011010001", b"10110000001101000100001010100000"), -- -6.55783e-10 + -5.1438e-39 = -6.55783e-10
	(b"10111111110000101011010101111100", b"00000000000000000000000000000000"),
	(b"10000000000100101100110110010001", b"10111111110000101011010101111100"), -- -1.52116 + -1.72678e-39 = -1.52116
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010011100111001110001000", b"10000000010011100111001110001000"), -- 0 + -7.20461e-39 = -7.20461e-39
	(b"11100000110001100101001000100010", b"00000000000000000000000000000000"),
	(b"10000000000110010001011000100111", b"11100000110001100101001000100010"), -- -1.14324e+20 + -2.30383e-39 = -1.14324e+20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010001100100101010100", b"10000000001010001100100101010100"), -- -0 + -3.74564e-39 = -3.74564e-39
	(b"11100001110111010001100110000100", b"00000000000000000000000000000000"),
	(b"00000000010100101100101011001111", b"11100001110111010001100110000100"), -- -5.09821e+20 + 7.60326e-39 = -5.09821e+20
	(b"01001000110110110010001010010000", b"00000000000000000000000000000000"),
	(b"00000000010100010011111101111101", b"01001000110110110010001010010000"), -- 448788 + 7.46145e-39 = 448788
	(b"11001010001011010010101010101111", b"00000000000000000000000000000000"),
	(b"10000000001011110100001110011001", b"11001010001011010010101010101111"), -- -2.83716e+06 + -4.34052e-39 = -2.83716e+06
	(b"01011101110000110100000011111000", b"00000000000000000000000000000000"),
	(b"00000000010000000010000011000010", b"01011101110000110100000011111000"), -- 1.75869e+18 + 5.88922e-39 = 1.75869e+18
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000111000000010010110", b"00000000001000111000000010010110"), -- 0 + 3.26037e-39 = 3.26037e-39
	(b"00101001011011101100011101001010", b"00000000000000000000000000000000"),
	(b"10000000011010011101010110001011", b"00101001011011101100011101001010"), -- 5.30195e-14 + -9.71933e-39 = 5.30195e-14
	(b"11110101000001101000111001001111", b"00000000000000000000000000000000"),
	(b"00000000010110010101100100100111", b"11110101000001101000111001001111"), -- -1.7057e+32 + 8.20534e-39 = -1.7057e+32
	(b"01001001100101100110001001111010", b"00000000000000000000000000000000"),
	(b"10000000011100011111011000101001", b"01001001100101100110001001111010"), -- 1.23195e+06 + -1.04657e-38 = 1.23195e+06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000010110001001010101", b"10000000000000010110001001010101"), -- 0 + -1.2711e-40 = -1.2711e-40
	(b"01001100001010001100101011101000", b"00000000000000000000000000000000"),
	(b"10000000010001010000100101010010", b"01001100001010001100101011101000"), -- 4.4248e+07 + -6.33999e-39 = 4.4248e+07
	(b"11101000001000001000111011100101", b"00000000000000000000000000000000"),
	(b"00000000000101011010110101010000", b"11101000001000001000111011100101"), -- -3.03286e+24 + 1.99072e-39 = -3.03286e+24
	(b"00100000011111011010010100011000", b"00000000000000000000000000000000"),
	(b"00000000001001001110111011010000", b"00100000011111011010010100011000"), -- 2.14846e-19 + 3.39175e-39 = 2.14846e-19
	(b"10000110100011011110001110010101", b"00000000000000000000000000000000"),
	(b"10000000010000011001010010110000", b"10000110100011011110011110101110"), -- -5.33727e-35 + -6.02265e-39 = -5.33787e-35
	(b"01011011010010101000101101011100", b"00000000000000000000000000000000"),
	(b"00000000011001110101100101010111", b"01011011010010101000101101011100"), -- 5.70112e+16 + 9.49111e-39 = 5.70112e+16
	(b"00000011011100011000111000101000", b"00000000000000000000000000000000"),
	(b"00000000000010000110001100011010", b"00000011011100011101000101000001"), -- 7.09867e-37 + 7.70235e-40 = 7.10637e-37
	(b"11010010100010010101010010000011", b"00000000000000000000000000000000"),
	(b"10000000011111000101011101101011", b"11010010100010010101010010000011"), -- -2.94914e+11 + -1.1419e-38 = -2.94914e+11
	(b"11011000010001011100001001010001", b"00000000000000000000000000000000"),
	(b"00000000000011100101011001010100", b"11011000010001011100001001010001"), -- -8.69753e+14 + 1.31667e-39 = -8.69753e+14
	(b"11000100010010101111101111101100", b"00000000000000000000000000000000"),
	(b"00000000001111110110100110110011", b"11000100010010101111101111101100"), -- -811.936 + 5.82355e-39 = -811.936
	(b"00101010000010101111011110111000", b"00000000000000000000000000000000"),
	(b"00000000011110110101010100010000", b"00101010000010101111011110111000"), -- 1.23428e-13 + 1.13263e-38 = 1.23428e-13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010010111010110100001000", b"11111111100000000000000000000000"), -- -inf + 6.94973e-39 = -inf
	(b"00110111001101110000100000010100", b"00000000000000000000000000000000"),
	(b"10000000011010100000000100011111", b"00110111001101110000100000010100"), -- 1.09095e-05 + -9.73496e-39 = 1.09095e-05
	(b"10111100100010011000110101000000", b"00000000000000000000000000000000"),
	(b"10000000000110010101111111011000", b"10111100100010011000110101000000"), -- -0.016791 + -2.33027e-39 = -0.016791
	(b"01001010100100100000010100101101", b"00000000000000000000000000000000"),
	(b"10000000000111011011110010011100", b"01001010100100100000010100101101"), -- 4.78479e+06 + -2.73089e-39 = 4.78479e+06
	(b"11100010010010101100010001001110", b"00000000000000000000000000000000"),
	(b"10000000011010101000011001010110", b"11100010010010101100010001001110"), -- -9.35097e+20 + -9.78275e-39 = -9.35097e+20
	(b"11001111000000001111001110000011", b"00000000000000000000000000000000"),
	(b"00000000000001011101110100000111", b"11001111000000001111001110000011"), -- -2.16344e+09 + 5.38467e-40 = -2.16344e+09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000110110000111100001000", b"01111111100000000000000000000000"), -- inf + 2.48495e-39 = inf
	(b"01000101111000001111000100110100", b"00000000000000000000000000000000"),
	(b"10000000010101001110010010010001", b"01000101111000001111000100110100"), -- 7198.15 + -7.79618e-39 = 7198.15
	(b"01000010010000011100000100010011", b"00000000000000000000000000000000"),
	(b"00000000010100100111010110101001", b"01000010010000011100000100010011"), -- 48.4385 + 7.57272e-39 = 48.4385
	(b"10000000000000000000000000010101", b"00000000000000000000000000000000"),
	(b"10000000000100010001000011101000", b"10000000000100010001000011111101"), -- -2.94273e-44 + -1.56727e-39 = -1.5673e-39
	(b"10101000101100001010001000000110", b"00000000000000000000000000000000"),
	(b"00000000011000001101110000011101", b"10101000101100001010001000000110"), -- -1.96102e-14 + 8.89517e-39 = -1.96102e-14
	(b"01110010000110100010000111111101", b"00000000000000000000000000000000"),
	(b"00000000000001010110110010111001", b"01110010000110100010000111111101"), -- 3.05291e+30 + 4.9818e-40 = 3.05291e+30
	(b"00010101101000010011011001011000", b"00000000000000000000000000000000"),
	(b"00000000010101100100110100000011", b"00010101101000010011011001011000"), -- 6.51131e-26 + 7.92548e-39 = 6.51131e-26
	(b"11011011000100111100111010111000", b"00000000000000000000000000000000"),
	(b"00000000010000000001111010100101", b"11011011000100111100111010111000"), -- -4.16041e+16 + 5.88846e-39 = -4.16041e+16
	(b"10011100010010010111010110100100", b"00000000000000000000000000000000"),
	(b"10000000011100011111100100010101", b"10011100010010010111010110100100"), -- -6.66574e-22 + -1.04668e-38 = -6.66574e-22
	(b"01010010101100011100000101011101", b"00000000000000000000000000000000"),
	(b"10000000010000111001000000100010", b"01010010101100011100000101011101"), -- 3.81727e+11 + -6.20468e-39 = 3.81727e+11
	(b"00011111010100111100101100000111", b"00000000000000000000000000000000"),
	(b"00000000000000101010110101011110", b"00011111010100111100101100000111"), -- 4.48489e-20 + 2.45863e-40 = 4.48489e-20
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011110011011101100110110", b"11111111100000000000000000000000"), -- -inf + 1.11793e-38 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000110011000100110011", b"01111111100000000000000000000000"), -- inf + 2.93156e-40 = inf
	(b"00010101111001011100010010001111", b"00000000000000000000000000000000"),
	(b"10000000010100111001111100001100", b"00010101111001011100010010001111"), -- 9.28025e-26 + -7.6794e-39 = 9.28025e-26
	(b"11110011101100100110010101010001", b"00000000000000000000000000000000"),
	(b"10000000010110011111001011001000", b"11110011101100100110010101010001"), -- -2.82679e+31 + -8.26045e-39 = -2.82679e+31
	(b"01110011101010101110110011011111", b"00000000000000000000000000000000"),
	(b"00000000010110100111011000011100", b"01110011101010101110110011011111"), -- 2.70842e+31 + 8.30756e-39 = 2.70842e+31
	(b"00111011111010001010110000011110", b"00000000000000000000000000000000"),
	(b"00000000011011010111110001101101", b"00111011111010001010110000011110"), -- 0.0071006 + 1.00547e-38 = 0.0071006
	(b"01111101110110001000101011001101", b"00000000000000000000000000000000"),
	(b"00000000010010001101010000100010", b"01111101110110001000101011001101"), -- 3.59792e+37 + 6.68825e-39 = 3.59792e+37
	(b"10001000111000000000110010001000", b"00000000000000000000000000000000"),
	(b"00000000010110111011101010110101", b"10001000111000000000110000101100"), -- -1.34845e-33 + 8.42401e-39 = -1.34844e-33
	(b"10011111011010001110000110000001", b"00000000000000000000000000000000"),
	(b"00000000000010100010101111010110", b"10011111011010001110000110000001"), -- -4.93144e-20 + 9.3408e-40 = -4.93144e-20
	(b"01011001000111001010110101110011", b"00000000000000000000000000000000"),
	(b"10000000001110011101111100010010", b"01011001000111001010110101110011"), -- 2.7563e+15 + -5.31465e-39 = 2.7563e+15
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001010101100110010111", b"11111111100000000000000000000000"), -- -inf + 9.30752e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001101100000101000010011", b"01111111100000000000000000000000"), -- inf + 4.96273e-39 = inf
	(b"10010111001011000010011110110000", b"00000000000000000000000000000000"),
	(b"00000000011110011111110010011110", b"10010111001011000010011110110000"), -- -5.56263e-25 + 1.12027e-38 = -5.56263e-25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010010011100110111011001", b"11111111100000000000000000000000"), -- -inf + -6.77784e-39 = -inf
	(b"01101101100110010110100010010110", b"00000000000000000000000000000000"),
	(b"10000000010001010111110010110110", b"01101101100110010110100010010110"), -- 5.93471e+27 + -6.38139e-39 = 5.93471e+27
	(b"00110001101110000010010110010001", b"00000000000000000000000000000000"),
	(b"10000000010101110110001000100000", b"00110001101110000010010110010001"), -- 5.35938e-09 + -8.02489e-39 = 5.35938e-09
	(b"00011010000111000001111000110111", b"00000000000000000000000000000000"),
	(b"00000000000011110100000011010001", b"00011010000111000001111000110111"), -- 3.22845e-23 + 1.40078e-39 = 3.22845e-23
	(b"00110000011010001110101110110000", b"00000000000000000000000000000000"),
	(b"10000000011100111100101001010011", b"00110000011010001110101110110000"), -- 8.4736e-10 + -1.06337e-38 = 8.4736e-10
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101011000011110001101", b"10000000011101011000011110001101"), -- -0 + -1.07934e-38 = -1.07934e-38
	(b"01101100000100100101100001010010", b"00000000000000000000000000000000"),
	(b"00000000000011100011010011001111", b"01101100000100100101100001010010"), -- 7.07681e+26 + 1.30464e-39 = 7.07681e+26
	(b"00000011010011111011111110000100", b"00000000000000000000000000000000"),
	(b"10000000000010100100110011110000", b"00000011010011110110110100011100"), -- 6.10517e-37 + -9.45955e-40 = 6.09571e-37
	(b"00010101110111001111110010010010", b"00000000000000000000000000000000"),
	(b"00000000000001111100010100100010", b"00010101110111001111110010010010"), -- 8.92558e-26 + 7.13566e-40 = 8.92558e-26
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010100111100001000010011", b"00000000010100111100001000010011"), -- 0 + 7.69197e-39 = 7.69197e-39
	(b"11001001011100000010000100010111", b"00000000000000000000000000000000"),
	(b"00000000000001000001000011101100", b"11001001011100000010000100010111"), -- -983569 + 3.73412e-40 = -983569
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110000000001111101011", b"10000000001110000000001111101011"), -- 0 + -5.14419e-39 = -5.14419e-39
	(b"11010011001010101110000011010100", b"00000000000000000000000000000000"),
	(b"10000000001110001100110101110011", b"11010011001010101110000011010100"), -- -7.33916e+11 + -5.21649e-39 = -7.33916e+11
	(b"11011010101001100100111000011111", b"00000000000000000000000000000000"),
	(b"00000000001100010000111000011010", b"11011010101001100100111000011111"), -- -2.34054e+16 + 4.505e-39 = -2.34054e+16
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010000100001001011111", b"10000000001010000100001001011111"), -- -0 + -3.69723e-39 = -3.69723e-39
	(b"11111011000001110001010000000010", b"00000000000000000000000000000000"),
	(b"00000000011100100111100110011011", b"11111011000001110001010000000010"), -- -7.01366e+35 + 1.05129e-38 = -7.01366e+35
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001011111001010011010", b"01111111100000000000000000000000"), -- inf + 6.42368e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111011111110101100001", b"11111111100000000000000000000000"), -- -inf + 2.75412e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001000101011101110101011", b"11111111100000000000000000000000"), -- -inf + -3.18973e-39 = -inf
	(b"01100110100110110110110101100111", b"00000000000000000000000000000000"),
	(b"00000000011000111011100001001010", b"01100110100110110110110101100111"), -- 3.66992e+23 + 9.15782e-39 = 3.66992e+23
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010011001111001010111010", b"11111111100000000000000000000000"), -- -inf + -7.06657e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001101011111010000100", b"01111111100000000000000000000000"), -- inf + 9.43556e-39 = inf
	(b"00000000000000000000110100010100", b"00000000000000000000000000000000"),
	(b"10000000001110110100101001110011", b"10000000001110110011110101011111"), -- 4.69155e-42 + -5.445e-39 = -5.44031e-39
	(b"11101101000101011001100110101110", b"00000000000000000000000000000000"),
	(b"00000000001010011001000001101010", b"11101101000101011001100110101110"), -- -2.89369e+27 + 3.81706e-39 = -2.89369e+27
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010111111100010111111101", b"01111111100000000000000000000000"), -- inf + 8.7954e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011111100010110000000111", b"11111111100000000000000000000000"), -- -inf + 1.15871e-38 = -inf
	(b"10001111111111110001100011001110", b"00000000000000000000000000000000"),
	(b"10000000011001101100011011001100", b"10001111111111110001100011001110"), -- -2.51545e-29 + -9.43854e-39 = -2.51545e-29
	(b"00000000000011000100011000000111", b"00000000000000000000000000000000"),
	(b"10000000000000100011010001100100", b"00000000000010100001000110100011"), -- 1.12715e-39 + -2.02465e-40 = 9.24682e-40
	(b"01111001100010010011001101011111", b"00000000000000000000000000000000"),
	(b"00000000010011110011100110010010", b"01111001100010010011001101011111"), -- 8.90483e+34 + 7.27566e-39 = 8.90483e+34
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111100100100101110111", b"11111111100000000000000000000000"), -- -inf + -8.65889e-39 = -inf
	(b"10110101110111010001100010110010", b"00000000000000000000000000000000"),
	(b"00000000000000100010111010110000", b"10110101110111010001100010110010"), -- -1.6473e-06 + 2.00419e-40 = -1.6473e-06
	(b"11000001110001111001110011011000", b"00000000000000000000000000000000"),
	(b"10000000010001100010110010011100", b"11000001110001111001110011011000"), -- -24.9516 + -6.44449e-39 = -24.9516
	(b"00000000001101111000110111110001", b"00000000000000000000000000000000"),
	(b"00000000001110000110111100011100", b"00000000011011111111110100001101"), -- 5.10187e-39 + 5.18265e-39 = 1.02845e-38
	(b"11110111111101100101011011001100", b"00000000000000000000000000000000"),
	(b"10000000000110010101000111001011", b"11110111111101100101011011001100"), -- -9.9927e+33 + -2.32523e-39 = -9.9927e+33
	(b"10101011000111110101010001011001", b"00000000000000000000000000000000"),
	(b"00000000000110101000011101000011", b"10101011000111110101010001011001"), -- -5.66052e-13 + 2.43625e-39 = -5.66052e-13
	(b"01000011110001111110110111011110", b"00000000000000000000000000000000"),
	(b"00000000011110000100101010001110", b"01000011110001111110110111011110"), -- 399.858 + 1.1047e-38 = 399.858
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000101111110011010101111", b"11111111100000000000000000000000"), -- -inf + 2.19497e-39 = -inf
	(b"10101110001100100001000000001010", b"00000000000000000000000000000000"),
	(b"10000000000000010110010101110010", b"10101110001100100001000000001010"), -- -4.04868e-11 + -1.28227e-40 = -4.04868e-11
	(b"01011001011110101000100111000011", b"00000000000000000000000000000000"),
	(b"10000000010101001001111111100011", b"01011001011110101000100111000011"), -- 4.40751e+15 + -7.77154e-39 = 4.40751e+15
	(b"11011110110011000001011101011000", b"00000000000000000000000000000000"),
	(b"00000000001010101000011011110001", b"11011110110011000001011101011000"), -- -7.35316e+18 + 3.9055e-39 = -7.35316e+18
	(b"00010110010000000101001000101010", b"00000000000000000000000000000000"),
	(b"10000000011001010011101110010111", b"00010110010000000101001000101010"), -- 1.55356e-25 + -9.29676e-39 = 1.55356e-25
	(b"01110111011011110001010100111110", b"00000000000000000000000000000000"),
	(b"10000000000000110011111011010011", b"01110111011011110001010100111110"), -- 4.84918e+33 + -2.98044e-40 = 4.84918e+33
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110001111111110010010", b"00000000010110001111111110010010"), -- -0 + 8.17321e-39 = 8.17321e-39
	(b"11010100011101110010001001001101", b"00000000000000000000000000000000"),
	(b"00000000011000110001100011001111", b"11010100011101110010001001001101"), -- -4.24573e+12 + 9.10061e-39 = -4.24573e+12
	(b"11100010000101010111010001111011", b"00000000000000000000000000000000"),
	(b"10000000010001100111111011111110", b"11100010000101010111010001111011"), -- -6.8924e+20 + -6.47404e-39 = -6.8924e+20
	(b"00110110100011001011111000010111", b"00000000000000000000000000000000"),
	(b"00000000010100101111010000001000", b"00110110100011001011111000010111"), -- 4.19445e-06 + 7.61805e-39 = 4.19445e-06
	(b"01111100100111110110011101000000", b"00000000000000000000000000000000"),
	(b"10000000010000110011110100011000", b"01111100100111110110011101000000"), -- 6.62135e+36 + -6.17489e-39 = 6.62135e+36
	(b"01010000000001000100100101111111", b"00000000000000000000000000000000"),
	(b"10000000010110101111011100010111", b"01010000000001000100100101111111"), -- 8.87764e+09 + -8.35383e-39 = 8.87764e+09
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011010111111101110011100", b"10000000011010111111101110011100"), -- 0 + -9.91666e-39 = -9.91666e-39
	(b"00101011100010010010100100011101", b"00000000000000000000000000000000"),
	(b"10000000011010000010011010011111", b"00101011100010010010100100011101"), -- 9.74585e-13 + -9.56475e-39 = 9.74585e-13
	(b"00101010100100011001110000000011", b"00000000000000000000000000000000"),
	(b"00000000001001001111111110000011", b"00101010100100011001110000000011"), -- 2.58654e-13 + 3.39774e-39 = 2.58654e-13
	(b"11110100111001110101111100111001", b"00000000000000000000000000000000"),
	(b"10000000000010010001000001010000", b"11110100111001110101111100111001"), -- -1.46649e+32 + -8.32371e-40 = -1.46649e+32
	(b"11001110100101010100101101011100", b"00000000000000000000000000000000"),
	(b"10000000000100010000001010101001", b"11001110100101010100101101011100"), -- -1.25237e+09 + -1.56216e-39 = -1.25237e+09
	(b"11010001010100001000000010011110", b"00000000000000000000000000000000"),
	(b"10000000001110011000100100100100", b"11010001010100001000000010011110"), -- -5.59694e+10 + -5.28382e-39 = -5.59694e+10
	(b"11001010000110101101000100000010", b"00000000000000000000000000000000"),
	(b"00000000010000101001011110000100", b"11001010000110101101000100000010"), -- -2.53651e+06 + 6.1155e-39 = -2.53651e+06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000001001110100000110", b"10000000011000001001110100000110"), -- -0 + -8.87254e-39 = -8.87254e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011000011101100001110111", b"11111111100000000000000000000000"), -- -inf + 8.9857e-39 = -inf
	(b"11101011000001001010100111101010", b"00000000000000000000000000000000"),
	(b"00000000010110001111111101010001", b"11101011000001001010100111101010"), -- -1.60381e+26 + 8.17311e-39 = -1.60381e+26
	(b"01001110111111011000001110110101", b"00000000000000000000000000000000"),
	(b"10000000000100001010010111010001", b"01001110111111011000001110110101"), -- 2.12663e+09 + -1.52885e-39 = 2.12663e+09
	(b"01101101000111011100110000100010", b"00000000000000000000000000000000"),
	(b"00000000011011011110010110011000", b"01101101000111011100110000100010"), -- 3.05225e+27 + 1.00924e-38 = 3.05225e+27
	(b"00010111110001101110101010000111", b"00000000000000000000000000000000"),
	(b"00000000011010001000110011000011", b"00010111110001101110101010000111"), -- 1.28547e-24 + 9.60139e-39 = 1.28547e-24
	(b"10011101111011001010111000011100", b"00000000000000000000000000000000"),
	(b"00000000000101111001011001101000", b"10011101111011001010111000011100"), -- -6.26487e-21 + 2.16617e-39 = -6.26487e-21
	(b"11101010001110010011000000001101", b"00000000000000000000000000000000"),
	(b"10000000010110011000111101011111", b"11101010001110010011000000001101"), -- -5.59695e+25 + -8.22479e-39 = -5.59695e+25
	(b"01100110111101010111101100111101", b"00000000000000000000000000000000"),
	(b"10000000011111110100000000010001", b"01100110111101010111101100111101"), -- 5.79627e+23 + -1.16861e-38 = 5.79627e+23
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000010001100100010011", b"01111111100000000000000000000000"), -- inf + -1.0083e-40 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000001111100001000101", b"01111111100000000000000000000000"), -- inf + 8.90623e-41 = inf
	(b"11010011110110011011001110100100", b"00000000000000000000000000000000"),
	(b"10000000000011001011010100010111", b"11010011110110011011001110100100"), -- -1.87004e+12 + -1.16699e-39 = -1.87004e+12
	(b"10101101010101010001100110101101", b"00000000000000000000000000000000"),
	(b"00000000001000101010010101101000", b"10101101010101010001100110101101"), -- -1.21133e-11 + 3.18174e-39 = -1.21133e-11
	(b"10000000000000000000000100000011", b"00000000000000000000000000000000"),
	(b"10000000011110111001111110011001", b"10000000011110111010000010011100"), -- -3.62936e-43 + -1.1353e-38 = -1.13534e-38
	(b"00101101011010101010100010011010", b"00000000000000000000000000000000"),
	(b"10000000011110010001101001111100", b"00101101011010101010100010011010"), -- 1.33388e-11 + -1.11216e-38 = 1.33388e-11
	(b"10000000000000000000000000000110", b"00000000000000000000000000000000"),
	(b"00000000001000110101000011111101", b"00000000001000110101000011110111"), -- -8.40779e-45 + 3.2433e-39 = 3.24329e-39
	(b"11010110011011101111100110111111", b"00000000000000000000000000000000"),
	(b"00000000011010000101011111011010", b"11010110011011101111100110111111"), -- -6.56891e+13 + 9.58241e-39 = -6.56891e+13
	(b"01001010101001001010101110111000", b"00000000000000000000000000000000"),
	(b"10000000010011100110000001000010", b"01001010101001001010101110111000"), -- 5.39593e+06 + -7.1977e-39 = 5.39593e+06
	(b"00111110001100101011110101101010", b"00000000000000000000000000000000"),
	(b"10000000000101011010001000010111", b"00111110001100101011110101101010"), -- 0.174551 + -1.98669e-39 = 0.174551
	(b"11111110001100001101011101101111", b"00000000000000000000000000000000"),
	(b"10000000001111100100000011111000", b"11111110001100001101011101101111"), -- -5.87657e+37 + -5.71711e-39 = -5.87657e+37
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011010000000100011011111", b"11111111100000000000000000000000"), -- -inf + 9.55407e-39 = -inf
	(b"01000101000101110110101100000011", b"00000000000000000000000000000000"),
	(b"10000000010000110010100011011010", b"01000101000101110110101100000011"), -- 2422.69 + -6.16763e-39 = 2422.69
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000101010011001000011110", b"00000000000101010011001000011110"), -- -0 + 1.94652e-39 = 1.94652e-39
	(b"00001010101110000101000110101111", b"00000000000000000000000000000000"),
	(b"00000000001011100000100011101110", b"00001010101110000101000110110010"), -- 1.77493e-32 + 4.22764e-39 = 1.77493e-32
	(b"10110101101100000000011110010000", b"00000000000000000000000000000000"),
	(b"00000000001000011000000100011011", b"10110101101100000000011110010000"), -- -1.31152e-06 + 3.07689e-39 = -1.31152e-06
	(b"10111110100010000101000100010010", b"00000000000000000000000000000000"),
	(b"10000000011101101111010110011011", b"10111110100010000101000100010010"), -- -0.266244 + -1.09247e-38 = -0.266244
	(b"11000111000100101111000110001100", b"00000000000000000000000000000000"),
	(b"00000000010110110100100110101001", b"11000111000100101111000110001100"), -- -37617.5 + 8.38345e-39 = -37617.5
	(b"10001010000010011101101110111010", b"00000000000000000000000000000000"),
	(b"10000000010101101011100111001010", b"10001010000010011101101111000101"), -- -6.63764e-33 + -7.9645e-39 = -6.63764e-33
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100001111001110110011", b"01111111100000000000000000000000"), -- inf + -1.0373e-38 = inf
	(b"00000000000000000000000001001110", b"00000000000000000000000000000000"),
	(b"00000000010000011010000101101110", b"00000000010000011010000110111100"), -- 1.09301e-43 + 6.02722e-39 = 6.02733e-39
	(b"00111001101001100001000011101111", b"00000000000000000000000000000000"),
	(b"10000000001011101101110101010111", b"00111001101001100001000011101111"), -- 0.000316746 + -4.30383e-39 = 0.000316746
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001110001111011110001", b"00000000010001110001111011110001"), -- -0 + 6.53142e-39 = 6.53142e-39
	(b"00100001000010110010000000000011", b"00000000000000000000000000000000"),
	(b"10000000001110110111010011110000", b"00100001000010110010000000000011"), -- 4.71374e-19 + -5.46024e-39 = 4.71374e-19
	(b"01001000000111011110110100111100", b"00000000000000000000000000000000"),
	(b"10000000000110110101101000110000", b"01001000000111011110110100111100"), -- 161717 + -2.51191e-39 = 161717
	(b"11100110000001011001101110010100", b"00000000000000000000000000000000"),
	(b"00000000010010001110000010000010", b"11100110000001011001101110010100"), -- -1.57736e+23 + 6.69269e-39 = -1.57736e+23
	(b"10010010010111110100001010110001", b"00000000000000000000000000000000"),
	(b"10000000000011000101110110100101", b"10010010010111110100001010110001"), -- -7.04486e-28 + -1.13562e-39 = -7.04486e-28
	(b"01000001001000110001010011111000", b"00000000000000000000000000000000"),
	(b"00000000011111010001011100000011", b"01000001001000110001010011111000"), -- 10.1926 + 1.14877e-38 = 10.1926
	(b"00000000000000000000000001100101", b"00000000000000000000000000000000"),
	(b"10000000000111111000110001000111", b"10000000000111111000101111100010"), -- 1.41531e-43 + -2.89722e-39 = -2.89708e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000000111100010111010", b"00000000001000000111100010111010"), -- -0 + 2.98204e-39 = 2.98204e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110110100111011110001", b"10000000011110110100111011110001"), -- 0 + -1.13241e-38 = -1.13241e-38
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010100010011000001011100", b"00000000010100010011000001011100"), -- 0 + 7.45602e-39 = 7.45602e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010000101100100010000000", b"00000000010000101100100010000000"), -- -0 + 6.13307e-39 = 6.13307e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011101011010001011001", b"00000000000011101011010001011001"), -- -0 + 1.35039e-39 = 1.35039e-39
	(b"11011110100001010001101010111011", b"00000000000000000000000000000000"),
	(b"00000000001000100011001011010001", b"11011110100001010001101010111011"), -- -4.79559e+18 + 3.14064e-39 = -4.79559e+18
	(b"10100001101000010100000011100101", b"00000000000000000000000000000000"),
	(b"10000000001000001100010000111000", b"10100001101000010100000011100101"), -- -1.0927e-18 + -3.00913e-39 = -1.0927e-18
	(b"10100000010100001001100100011001", b"00000000000000000000000000000000"),
	(b"10000000000010011101111011011011", b"10100000010100001001100100011001"), -- -1.76689e-19 + -9.06465e-40 = -1.76689e-19
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000011100011010100100", b"10000000011000011100011010100100"), -- -0 + -8.9793e-39 = -8.9793e-39
	(b"01011001011111001110001100000100", b"00000000000000000000000000000000"),
	(b"00000000001111101000001001011110", b"01011001011111001110001100000100"), -- 4.44883e+15 + 5.74057e-39 = 4.44883e+15
	(b"11001010001001111101010010100101", b"00000000000000000000000000000000"),
	(b"00000000001111101010101000100111", b"11001010001001111101010010100101"), -- -2.74974e+06 + 5.75484e-39 = -2.74974e+06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001011000110000011010", b"10000000011001011000110000011010"), -- 0 + -9.32564e-39 = -9.32564e-39
	(b"01110011110110011110101110110010", b"00000000000000000000000000000000"),
	(b"00000000011010011001100100111111", b"01110011110110011110101110110010"), -- 3.45309e+31 + 9.6977e-39 = 3.45309e+31
	(b"00110010011001010010010011110000", b"00000000000000000000000000000000"),
	(b"10000000001100111100011000001100", b"00110010011001010010010011110000"), -- 1.3338e-08 + -4.75466e-39 = 1.3338e-08
	(b"10011101011000001000111011001001", b"00000000000000000000000000000000"),
	(b"00000000001000001111100101101100", b"10011101011000001000111011001001"), -- -2.972e-21 + 3.02821e-39 = -2.972e-21
	(b"10001010001011101001001011101111", b"00000000000000000000000000000000"),
	(b"10000000011011001110010011110010", b"10001010001011101001001011111101"), -- -8.40543e-33 + -1.00004e-38 = -8.40544e-33
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011111000111000111110010", b"00000000011111000111000111110010"), -- -0 + 1.14285e-38 = 1.14285e-38
	(b"11000001100111000001111010101110", b"00000000000000000000000000000000"),
	(b"00000000001110010100100010001001", b"11000001100111000001111010101110"), -- -19.515 + 5.26064e-39 = -19.515
	(b"11010100001101001100011110001110", b"00000000000000000000000000000000"),
	(b"10000000010100010010111001000010", b"11010100001101001100011110001110"), -- -3.10577e+12 + -7.45527e-39 = -3.10577e+12
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011010101010110111011101", b"00000000011010101010110111011101"), -- 0 + 9.79693e-39 = 9.79693e-39
	(b"01010100101110101010100000101110", b"00000000000000000000000000000000"),
	(b"00000000010000101111001100011101", b"01010100101110101010100000101110"), -- 6.41348e+12 + 6.14836e-39 = 6.41348e+12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110101100011010000010", b"11111111100000000000000000000000"), -- -inf + 5.39767e-39 = -inf
	(b"10100110110000101000101000011010", b"00000000000000000000000000000000"),
	(b"10000000010001001111001111001100", b"10100110110000101000101000011010"), -- -1.34989e-15 + -6.33227e-39 = -1.34989e-15
	(b"11100010001110111111000100011111", b"00000000000000000000000000000000"),
	(b"00000000000110011010100100011001", b"11100010001110111111000100011111"), -- -8.66729e+20 + 2.35655e-39 = -8.66729e+20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001110100011100001110", b"10000000001001110100011100001110"), -- -0 + -3.60707e-39 = -3.60707e-39
	(b"01100100111101111011110111010101", b"00000000000000000000000000000000"),
	(b"00000000000100101101101011000010", b"01100100111101111011110111010101"), -- 3.65602e+22 + 1.73151e-39 = 3.65602e+22
	(b"11111010010110100001111100001001", b"00000000000000000000000000000000"),
	(b"10000000010011011100101001101110", b"11111010010110100001111100001001"), -- -2.83138e+35 + -7.14395e-39 = -2.83138e+35
	(b"10110101101111001000001010110111", b"00000000000000000000000000000000"),
	(b"10000000010001000110001100010111", b"10110101101111001000001010110111"), -- -1.40451e-06 + -6.28036e-39 = -1.40451e-06
	(b"11001000001001010110000100011110", b"00000000000000000000000000000000"),
	(b"00000000000110110110010101111011", b"11001000001001010110000100011110"), -- -169348 + 2.51596e-39 = -169348
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001100011111111100110010", b"10000000001100011111111100110010"), -- 0 + -4.59149e-39 = -4.59149e-39
	(b"01111000001010110001010010111000", b"00000000000000000000000000000000"),
	(b"00000000000110100101100011011000", b"01111000001010110001010010111000"), -- 1.38797e+34 + 2.41959e-39 = 1.38797e+34
	(b"00011000011000111010010111011011", b"00000000000000000000000000000000"),
	(b"00000000011101001100000001100011", b"00011000011000111010010111011011"), -- 2.94228e-24 + 1.07219e-38 = 2.94228e-24
	(b"10110101010000101001111101010001", b"00000000000000000000000000000000"),
	(b"10000000011001010011100100001010", b"10110101010000101001111101010001"), -- -7.25025e-07 + -9.29585e-39 = -7.25025e-07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000110111000100101000", b"00000000001000110111000100101000"), -- -0 + 3.25484e-39 = 3.25484e-39
	(b"10110010011000000100100001100010", b"00000000000000000000000000000000"),
	(b"10000000010011111101010110000000", b"10110010011000000100100001100010"), -- -1.3055e-08 + -7.33159e-39 = -1.3055e-08
	(b"00111110100000010010100110010001", b"00000000000000000000000000000000"),
	(b"10000000011000001001110000111110", b"00111110100000010010100110010001"), -- 0.25227 + -8.87226e-39 = 0.25227
	(b"11000110000001011010011010101010", b"00000000000000000000000000000000"),
	(b"00000000011010111111110000011110", b"11000110000001011010011010101010"), -- -8553.67 + 9.91684e-39 = -8553.67
	(b"10101101000101000101011100100101", b"00000000000000000000000000000000"),
	(b"00000000011100101101010010000000", b"10101101000101000101011100100101"), -- -8.43218e-12 + 1.05455e-38 = -8.43218e-12
	(b"11101101100111011010100110010010", b"00000000000000000000000000000000"),
	(b"10000000000111010010100101000111", b"11101101100111011010100110010010"), -- -6.09927e+27 + -2.67804e-39 = -6.09927e+27
	(b"11100001100110010011100000111010", b"00000000000000000000000000000000"),
	(b"00000000001110101110110000010000", b"11100001100110010011100000111010"), -- -3.533e+20 + 5.41114e-39 = -3.533e+20
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000001101110101001010", b"11111111100000000000000000000000"), -- -inf + -7.93836e-41 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111000101111000001101", b"00000000000111000101111000001101"), -- 0 + 2.60513e-39 = 2.60513e-39
	(b"00110001110001101111000100001010", b"00000000000000000000000000000000"),
	(b"00000000010101100011011111000010", b"00110001110001101111000100001010"), -- 5.78996e-09 + 7.91785e-39 = 5.78996e-09
	(b"01100111000100100000000110100010", b"00000000000000000000000000000000"),
	(b"10000000001001010111100101010001", b"01100111000100100000000110100010"), -- 6.89496e+23 + -3.44143e-39 = 6.89496e+23
	(b"01000001000001111000110111101001", b"00000000000000000000000000000000"),
	(b"10000000000001101111111011001000", b"01000001000001111000110111101001"), -- 8.47215 + -6.42411e-40 = 8.47215
	(b"11111110100011011100101000011101", b"00000000000000000000000000000000"),
	(b"10000000000110111011000001100011", b"11111110100011011100101000011101"), -- -9.42353e+37 + -2.54283e-39 = -9.42353e+37
	(b"11000010000010111100101111111010", b"00000000000000000000000000000000"),
	(b"00000000010100000000010000111001", b"11000010000010111100101111111010"), -- -34.9492 + 7.34835e-39 = -34.9492
	(b"10110101010111111110001000110001", b"00000000000000000000000000000000"),
	(b"10000000011000011000001000011111", b"10110101010111111110001000110001"), -- -8.34031e-07 + -8.95472e-39 = -8.34031e-07
	(b"00000011110011111101010010001011", b"00000000000000000000000000000000"),
	(b"10000000000101110101010100101011", b"00000011110011110111011100110110"), -- 1.22152e-36 + -2.14277e-39 = 1.21937e-36
	(b"10100100111101001111111111000011", b"00000000000000000000000000000000"),
	(b"10000000000100101111111010111111", b"10100100111101001111111111000011"), -- -1.06251e-16 + -1.74442e-39 = -1.06251e-16
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011011010011111111110101", b"10000000011011010011111111110101"), -- -0 + -1.0033e-38 = -1.0033e-38
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000001011000001100011", b"00000000000000001011000001100011"), -- 0 + 6.32756e-41 = 6.32756e-41
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110011011000111111111", b"01111111100000000000000000000000"), -- inf + -1.11759e-38 = inf
	(b"11110001010011011100010000111110", b"00000000000000000000000000000000"),
	(b"00000000011111101111000100011101", b"11110001010011011100010000111110"), -- -1.01891e+30 + 1.16578e-38 = -1.01891e+30
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011100101101110111010", b"00000000000011100101101110111010"), -- -0 + 1.3186e-39 = 1.3186e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010001001011110111011100", b"01111111100000000000000000000000"), -- inf + -6.31292e-39 = inf
	(b"10000100000110011111000110011100", b"00000000000000000000000000000000"),
	(b"00000000001011111011001010011000", b"10000100000110011001001000110111"), -- -1.8096e-36 + 4.38034e-39 = -1.80522e-36
	(b"00001101000010000010100111101100", b"00000000000000000000000000000000"),
	(b"10000000001111110111101000010011", b"00001101000010000010100111101100"), -- 4.19587e-31 + -5.82943e-39 = 4.19587e-31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111111001000010111001", b"11111111100000000000000000000000"), -- -inf + 2.89882e-39 = -inf
	(b"00110100000011010011010001111000", b"00000000000000000000000000000000"),
	(b"00000000010110011100110010011101", b"00110100000011010011010001111000"), -- 1.31507e-07 + 8.24676e-39 = 1.31507e-07
	(b"00011110111110110000100001010110", b"00000000000000000000000000000000"),
	(b"10000000011000110111001001110101", b"00011110111110110000100001010110"), -- 2.65791e-20 + -9.13277e-39 = 2.65791e-20
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001101011110011111001", b"11111111100000000000000000000000"), -- -inf + -9.43501e-39 = -inf
	(b"11010101110010111010100011001011", b"00000000000000000000000000000000"),
	(b"00000000011111010111011001110011", b"11010101110010111010100011001011"), -- -2.79907e+13 + 1.15219e-38 = -2.79907e+13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010000011000101011100010", b"11111111100000000000000000000000"), -- -inf + -6.01913e-39 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000110010001101000101101", b"10000000000110010001101000101101"), -- 0 + -2.30528e-39 = -2.30528e-39
	(b"01000100010100000010110111001111", b"00000000000000000000000000000000"),
	(b"10000000001000101001011011010111", b"01000100010100000010110111001111"), -- 832.716 + -3.17652e-39 = 832.716
	(b"00101100010100101100001100010111", b"00000000000000000000000000000000"),
	(b"10000000000111001110010110000010", b"00101100010100101100001100010111"), -- 2.99511e-12 + -2.65373e-39 = 2.99511e-12
	(b"00000100001001011110011110111100", b"00000000000000000000000000000000"),
	(b"00000000011100011010101011111111", b"00000100001001101100101100010010"), -- 1.95021e-36 + 1.04388e-38 = 1.96065e-36
	(b"01001011100110000010001111011101", b"00000000000000000000000000000000"),
	(b"10000000000101001110000010111111", b"01001011100110000010001111011101"), -- 1.99413e+07 + -1.91733e-39 = 1.99413e+07
	(b"01111000101011111011001100101010", b"00000000000000000000000000000000"),
	(b"00000000011101000110011011010001", b"01111000101011111011001100101010"), -- 2.85089e+34 + 1.06898e-38 = 2.85089e+34
	(b"10000101100110001100110101100000", b"00000000000000000000000000000000"),
	(b"00000000010101010111001000011011", b"10000101100110001011100000000011"), -- -1.43695e-35 + 7.84695e-39 = -1.43616e-35
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011001110011100101011", b"01111111100000000000000000000000"), -- inf + 4.12369e-39 = inf
	(b"00001000000100111100110110010111", b"00000000000000000000000000000000"),
	(b"10000000001000101011011000001000", b"00001000000100111100110101010010"), -- 4.44779e-34 + -3.18771e-39 = 4.44776e-34
	(b"11011010001101110110100111110101", b"00000000000000000000000000000000"),
	(b"10000000000001111000111000000110", b"11011010001101110110100111110101"), -- -1.29066e+16 + -6.93797e-40 = -1.29066e+16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111100010010110000101", b"01111111100000000000000000000000"), -- inf + -8.646e-39 = inf
	(b"10101000010110110101010101111100", b"00000000000000000000000000000000"),
	(b"00000000010111100100011101001100", b"10101000010110110101010101111100"), -- -1.21755e-14 + 8.65811e-39 = -1.21755e-14
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011110101100111111111", b"01111111100000000000000000000000"), -- inf + -1.40982e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101011011011100110101", b"10000000011101011011011100110101"), -- 0 + -1.08105e-38 = -1.08105e-38
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110000100000000001110", b"00000000001110000100000000001110"), -- -0 + 5.16577e-39 = 5.16577e-39
	(b"11000010000001100110101110101001", b"00000000000000000000000000000000"),
	(b"10000000011101101100000101010010", b"11000010000001100110101110101001"), -- -33.6051 + -1.09059e-38 = -33.6051
	(b"00100000110000110111001110101000", b"00000000000000000000000000000000"),
	(b"10000000010110111001001011101011", b"00100000110000110111001110101000"), -- 3.31108e-19 + -8.40973e-39 = 3.31108e-19
	(b"01101111110000011110011011011100", b"00000000000000000000000000000000"),
	(b"10000000001011101011100011110010", b"01101111110000011110011011011100"), -- 1.20019e+29 + -4.29078e-39 = 1.20019e+29
	(b"11010101101000010101101000000111", b"00000000000000000000000000000000"),
	(b"00000000011000010010010011000010", b"11010101101000010101101000000111"), -- -2.2176e+13 + 8.92123e-39 = -2.2176e+13
	(b"01101110110010001000111111010001", b"00000000000000000000000000000000"),
	(b"10000000000110000111100100000010", b"01101110110010001000111111010001"), -- 3.10354e+28 + -2.24746e-39 = 3.10354e+28
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000101111111100111000", b"00000000000000101111111100111000"), -- 0 + 2.75226e-40 = 2.75226e-40
	(b"11000110001011011010100110010010", b"00000000000000000000000000000000"),
	(b"10000000001101001001101101110100", b"11000110001011011010100110010010"), -- -11114.4 + -4.83121e-39 = -11114.4
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000101000100001101100", b"01111111100000000000000000000000"), -- inf + -9.04882e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110101000100001001100", b"11111111100000000000000000000000"), -- -inf + -5.37535e-39 = -inf
	(b"10010010101001000111110011000111", b"00000000000000000000000000000000"),
	(b"00000000010110011100001111001101", b"10010010101001000111110011000111"), -- -1.03806e-27 + 8.2436e-39 = -1.03806e-27
	(b"11010100101011001000101011100101", b"00000000000000000000000000000000"),
	(b"10000000001010111100110000110101", b"11010100101011001000101011100101"), -- -5.92852e+12 + -4.02218e-39 = -5.92852e+12
	(b"11101101101111101000001100111010", b"00000000000000000000000000000000"),
	(b"00000000011111000010100000000000", b"11101101101111101000001100111010"), -- -7.3701e+27 + 1.1402e-38 = -7.3701e+27
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010011001001011100110101", b"01111111100000000000000000000000"), -- inf + -7.03374e-39 = inf
	(b"10000011100000000000001100011110", b"00000000000000000000000000000000"),
	(b"10000000000001100011110001111010", b"10000011100000000001110000010000"), -- -7.52388e-37 + -5.72708e-40 = -7.52961e-37
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001110000110101001110", b"11111111100000000000000000000000"), -- -inf + -9.46383e-39 = -inf
	(b"00011110110111001001010011101011", b"00000000000000000000000000000000"),
	(b"00000000001100011001101101101001", b"00011110110111001001010011101011"), -- 2.3355e-20 + 4.55569e-39 = 2.3355e-20
	(b"00100000101100101111101001011110", b"00000000000000000000000000000000"),
	(b"00000000011010110101111100110111", b"00100000101100101111101001011110"), -- 3.03201e-19 + 9.86055e-39 = 3.03201e-19
	(b"10001011110010101011001110100010", b"00000000000000000000000000000000"),
	(b"00000000001100000100101011001010", b"10001011110010101011001110100001"), -- -7.80779e-32 + 4.43493e-39 = -7.80778e-32
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011000011101011101101110", b"11111111100000000000000000000000"), -- -inf + 8.98532e-39 = -inf
	(b"00000000000000000100100110000010", b"00000000000000000000000000000000"),
	(b"00000000001011001000011000001100", b"00000000001011001100111110001110"), -- 2.63696e-41 + 4.08885e-39 = 4.11522e-39
	(b"10100010000100101111101010100111", b"00000000000000000000000000000000"),
	(b"10000000010111111110001011110100", b"10100010000100101111101010100111"), -- -1.99194e-18 + -8.80579e-39 = -1.99194e-18
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011111111011101001010", b"10000000000011111111011101001010"), -- -0 + -1.46624e-39 = -1.46624e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001000001110111000101001", b"10000000001000001110111000101001"), -- 0 + -3.02417e-39 = -3.02417e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011001011100001100001", b"01111111100000000000000000000000"), -- inf + 1.16817e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011101001010001111100000", b"01111111100000000000000000000000"), -- inf + -1.07117e-38 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011001011011110101110", b"00000000011011001011011110101110"), -- -0 + 9.98413e-39 = 9.98413e-39
	(b"11100101100010101101001001111010", b"00000000000000000000000000000000"),
	(b"10000000011001001111010010000000", b"11100101100010101101001001111010"), -- -8.19461e+22 + -9.27126e-39 = -8.19461e+22
	(b"10001001010011101111111000111001", b"00000000000000000000000000000000"),
	(b"00000000000000111111101101110000", b"10001001010011101111111000110111"), -- -2.49159e-33 + 3.65705e-40 = -2.49159e-33
	(b"00000000000000001101001100100111", b"00000000000000000000000000000000"),
	(b"00000000001101100110101011110010", b"00000000001101110011111000011001"), -- 7.57472e-41 + 4.99748e-39 = 5.07323e-39
	(b"01011001110000011111010110001000", b"00000000000000000000000000000000"),
	(b"10000000010001000110010111011010", b"01011001110000011111010110001000"), -- 6.82433e+15 + -6.28135e-39 = 6.82433e+15
	(b"10101111110000111100011010000101", b"00000000000000000000000000000000"),
	(b"00000000001111011111010011111101", b"10101111110000111100011010000101"), -- -3.56113e-10 + 5.68985e-39 = -3.56113e-10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001110111011100011001", b"11111111100000000000000000000000"), -- -inf + -9.50178e-39 = -inf
	(b"00000010101010000010001111000011", b"00000000000000000000000000000000"),
	(b"10000000001001001111000001111000", b"00000010101001011101010010111100"), -- 2.47059e-37 + -3.39234e-39 = 2.43667e-37
	(b"10101010001000000011100100110101", b"00000000000000000000000000000000"),
	(b"00000000010111010001110011111001", b"10101010001000000011100100110101"), -- -1.42307e-13 + 8.55109e-39 = -1.42307e-13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101011110010111010100", b"01111111100000000000000000000000"), -- inf + -4.94973e-39 = inf
	(b"00100000000101000011110001110110", b"00000000000000000000000000000000"),
	(b"00000000011101101001111010110111", b"00100000000101000011110001110110"), -- 1.25561e-19 + 1.08935e-38 = 1.25561e-19
	(b"10000101010010110011111000101001", b"00000000000000000000000000000000"),
	(b"00000000010011001011101000001010", b"10000101010010110001011111001100"), -- -9.55643e-36 + 7.04624e-39 = -9.54938e-36
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001100010010010101000000", b"11111111100000000000000000000000"), -- -inf + 4.5133e-39 = -inf
	(b"01001000100100011111101111001101", b"00000000000000000000000000000000"),
	(b"00000000010001011111101011000101", b"01001000100100011111101111001101"), -- 298974 + 6.42661e-39 = 298974
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011000101001001100110111", b"00000000011000101001001100110111"), -- -0 + 9.05269e-39 = 9.05269e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111000010011000010001", b"01111111100000000000000000000000"), -- inf + -8.46252e-39 = inf
	(b"00100101000001110001110011000101", b"00000000000000000000000000000000"),
	(b"00000000011110100100001100001100", b"00100101000001110001110011000101"), -- 1.17191e-16 + 1.1228e-38 = 1.17191e-16
	(b"00101001100000000110001110100110", b"00000000000000000000000000000000"),
	(b"10000000011111110011101101000001", b"00101001100000000110001110100110"), -- 5.70163e-14 + -1.16844e-38 = 5.70163e-14
	(b"00010101001110010100000001110011", b"00000000000000000000000000000000"),
	(b"10000000010011101100000111101011", b"00010101001110010100000001110011"), -- 3.74113e-26 + -7.23273e-39 = 3.74113e-26
	(b"10110110001111110001001100010100", b"00000000000000000000000000000000"),
	(b"10000000011000101000010110110110", b"10110110001111110001001100010100"), -- -2.84723e-06 + -9.04785e-39 = -2.84723e-06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000111010000011001110011", b"10000000000111010000011001110011"), -- 0 + -2.66554e-39 = -2.66554e-39
	(b"11100000110110100100110001110010", b"00000000000000000000000000000000"),
	(b"10000000001000110001111101010001", b"11100000110110100100110001110010"), -- -1.25841e+20 + -3.22548e-39 = -1.25841e+20
	(b"10010010111100111101010111111111", b"00000000000000000000000000000000"),
	(b"10000000000100010100000111001101", b"10010010111100111101010111111111"), -- -1.53882e-27 + -1.58481e-39 = -1.53882e-27
	(b"10010010011011000100110100000101", b"00000000000000000000000000000000"),
	(b"00000000011110010100101010101001", b"10010010011011000100110100000101"), -- -7.45634e-28 + 1.11389e-38 = -7.45634e-28
	(b"00010111100100101001001010010011", b"00000000000000000000000000000000"),
	(b"10000000011010001110000000010101", b"00010111100100101001001010010011"), -- 9.47203e-25 + -9.63128e-39 = 9.47203e-25
	(b"10000000000000000001010001100000", b"00000000000000000000000000000000"),
	(b"10000000001011001111000011001101", b"10000000001011010000010100101101"), -- -7.30917e-42 + -4.12714e-39 = -4.13445e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010100001110101110111101", b"01111111100000000000000000000000"), -- inf + -7.43141e-39 = inf
	(b"11101000111000011100001111010010", b"00000000000000000000000000000000"),
	(b"10000000011010001000111001010011", b"11101000111000011100001111010010"), -- -8.52916e+24 + -9.60195e-39 = -8.52916e+24
	(b"01110001011010001100111011111110", b"00000000000000000000000000000000"),
	(b"00000000001101111111000110110100", b"01110001011010001100111011111110"), -- 1.15281e+30 + 5.13766e-39 = 1.15281e+30
	(b"00110000101011000000110001110001", b"00000000000000000000000000000000"),
	(b"10000000011100100011010011100100", b"00110000101011000000110001110001"), -- 1.25182e-09 + -1.04882e-38 = 1.25182e-09
	(b"11001011010001111001101000001000", b"00000000000000000000000000000000"),
	(b"00000000010001100111000110111101", b"11001011010001111001101000001000"), -- -1.30811e+07 + 6.46929e-39 = -1.30811e+07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001101001101011010100", b"11111111100000000000000000000000"), -- -inf + 6.06555e-40 = -inf
	(b"11010111000110000010100010000111", b"00000000000000000000000000000000"),
	(b"10000000010001010100000101000011", b"11010111000110000010100010000111"), -- -1.673e+14 + -6.36006e-39 = -1.673e+14
	(b"01110110110111001000100110111101", b"00000000000000000000000000000000"),
	(b"10000000000111111110111111000010", b"01110110110111001000100110111101"), -- 2.23652e+33 + -2.93291e-39 = 2.23652e+33
	(b"11101010000001100010101011000000", b"00000000000000000000000000000000"),
	(b"00000000001001010101000001111001", b"11101010000001100010101011000000"), -- -4.05495e+25 + 3.42678e-39 = -4.05495e+25
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010011111101100001111110", b"00000000010011111101100001111110"), -- 0 + 7.33267e-39 = 7.33267e-39
	(b"00101110001001101000100001011100", b"00000000000000000000000000000000"),
	(b"10000000010000001100101010111000", b"00101110001001101000100001011100"), -- 3.78651e-11 + -5.95019e-39 = 3.78651e-11
	(b"11011001110111001001100100110000", b"00000000000000000000000000000000"),
	(b"00000000000101100011111100001000", b"11011001110111001001100100110000"), -- -7.76162e+15 + 2.04299e-39 = -7.76162e+15
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001101110111100100011101", b"00000000001101110111100100011101"), -- -0 + 5.0944e-39 = 5.0944e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001001011111000001100000", b"00000000001001011111000001100000"), -- -0 + 3.48414e-39 = 3.48414e-39
	(b"01100010110101110000010100000011", b"00000000000000000000000000000000"),
	(b"00000000001110100111110010101011", b"01100010110101110000010100000011"), -- 1.98321e+21 + 5.37118e-39 = 1.98321e+21
	(b"00101100100001010010101001100100", b"00000000000000000000000000000000"),
	(b"10000000001111011011110001001011", b"00101100100001010010101001100100"), -- 3.78479e-12 + -5.66951e-39 = 3.78479e-12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010010000000001010001101", b"11111111100000000000000000000000"), -- -inf + 6.61307e-39 = -inf
	(b"10100000101100010010000000001000", b"00000000000000000000000000000000"),
	(b"00000000011100011000011000010010", b"10100000101100010010000000001000"), -- -3.00062e-19 + 1.04255e-38 = -3.00062e-19
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110110111101110101110", b"01111111100000000000000000000000"), -- inf + 5.46266e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011000111110111011101", b"01111111100000000000000000000000"), -- inf + 1.14718e-39 = inf
	(b"01101100000011101010100000101101", b"00000000000000000000000000000000"),
	(b"00000000010000011111000010110110", b"01101100000011101010100000101101"), -- 6.89847e+26 + 6.05566e-39 = 6.89847e+26
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011100011100110000010011", b"00000000011100011100110000010011"), -- 0 + 1.04506e-38 = 1.04506e-38
	(b"10111010011010100001000100011111", b"00000000000000000000000000000000"),
	(b"10000000011011111110100101101010", b"10111010011010100001000100011111"), -- -0.000892894 + -1.02775e-38 = -0.000892894
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001100100010001000111", b"11111111100000000000000000000000"), -- -inf + -3.51424e-39 = -inf
	(b"11001000000010101100000111000000", b"00000000000000000000000000000000"),
	(b"10000000011010101010110111010111", b"11001000000010101100000111000000"), -- -142087 + -9.79692e-39 = -142087
	(b"01000010101001011101000000110010", b"00000000000000000000000000000000"),
	(b"10000000001001110110011011111100", b"01000010101001011101000000110010"), -- 82.9066 + -3.61853e-39 = 82.9066
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001000101101011100011", b"10000000001001000101101011100011"), -- -0 + -3.33868e-39 = -3.33868e-39
	(b"00011110101101011110010001010010", b"00000000000000000000000000000000"),
	(b"00000000000001000011111001001110", b"00011110101101011110010001010010"), -- 1.92586e-20 + 3.89693e-40 = 1.92586e-20
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101010100011011110101", b"00000000011101010100011011110101"), -- 0 + 1.07702e-38 = 1.07702e-38
	(b"10001101000000111011100111011001", b"00000000000000000000000000000000"),
	(b"00000000011001101100101011101011", b"10001101000000111011100111011001"), -- -4.05912e-31 + 9.44001e-39 = -4.05912e-31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000011111000100100011", b"11111111100000000000000000000000"), -- -inf + -8.99455e-39 = -inf
	(b"10001001100101001110011110100101", b"00000000000000000000000000000000"),
	(b"00000000011110001000001001011000", b"10001001100101001110011110000111"), -- -3.58475e-33 + 1.1067e-38 = -3.58474e-33
	(b"00111100011111011000010100000000", b"00000000000000000000000000000000"),
	(b"00000000000101000010011000010001", b"00111100011111011000010100000000"), -- 0.0154736 + 1.85037e-39 = 0.0154736
	(b"00101001001110100001111010101101", b"00000000000000000000000000000000"),
	(b"00000000000111010101111101001000", b"00101001001110100001111010101101"), -- 4.13269e-14 + 2.69741e-39 = 4.13269e-14
	(b"01100011000001100001111111000111", b"00000000000000000000000000000000"),
	(b"10000000000000111010101010111000", b"01100011000001100001111111000111"), -- 2.47415e+21 + -3.36749e-40 = 2.47415e+21
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100101000110101010010", b"01111111100000000000000000000000"), -- inf + -1.70374e-39 = inf
	(b"01110110001001011110000110101101", b"00000000000000000000000000000000"),
	(b"10000000011110010110011110010101", b"01110110001001011110000110101101"), -- 8.41119e+32 + -1.11493e-38 = 8.41119e+32
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010101011110011011001", b"00000000001010101011110011011001"), -- 0 + 3.92484e-39 = 3.92484e-39
	(b"10001000110101001000000111110000", b"00000000000000000000000000000000"),
	(b"10000000001111101101100101101011", b"10001000110101001000001000101111"), -- -1.27898e-33 + -5.7718e-39 = -1.27899e-33
	(b"01010100100101111101011010100101", b"00000000000000000000000000000000"),
	(b"00000000010000100100101011001001", b"01010100100101111101011010100101"), -- 5.21713e+12 + 6.08797e-39 = 5.21713e+12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011100100001111000101", b"11111111100000000000000000000000"), -- -inf + 1.31001e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110101010111010111111", b"11111111100000000000000000000000"), -- -inf + 8.32788e-39 = -inf
	(b"10101001001110010100100011110101", b"00000000000000000000000000000000"),
	(b"00000000001010001101111100001000", b"10101001001110010100100011110101"), -- -4.11415e-14 + 3.75343e-39 = -4.11415e-14
	(b"00111111100101111011011100000101", b"00000000000000000000000000000000"),
	(b"10000000010011111100000111010111", b"00111111100101111011011100000101"), -- 1.18527 + -7.32454e-39 = 1.18527
	(b"10000010101011000010101010011011", b"00000000000000000000000000000000"),
	(b"00000000000000001000000110010110", b"10000010101011000010001010000010"), -- -2.52976e-37 + 4.64867e-41 = -2.52929e-37
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001111000000100001010111", b"10000000001111000000100001010111"), -- 0 + -5.51312e-39 = -5.51312e-39
	(b"01101010111010100100010111100111", b"00000000000000000000000000000000"),
	(b"10000000010011010010000111011111", b"01101010111010100100010111100111"), -- 1.41609e+26 + -7.08348e-39 = 1.41609e+26
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111001110000110011011", b"01111111100000000000000000000000"), -- inf + 2.65233e-39 = inf
	(b"11100001000111001001011011010000", b"00000000000000000000000000000000"),
	(b"10000000000010001101111111111100", b"11100001000111001001011011010000"), -- -1.80535e+20 + -8.15034e-40 = -1.80535e+20
	(b"11111110111110011111010100101000", b"00000000000000000000000000000000"),
	(b"00000000001010111011111101000000", b"11111110111110011111010100101000"), -- -1.66125e+38 + 4.01753e-39 = -1.66125e+38
	(b"11010100000010010001111000000101", b"00000000000000000000000000000000"),
	(b"10000000011010111001100000110101", b"11010100000010010001111000000101"), -- -2.35566e+12 + -9.881e-39 = -2.35566e+12
	(b"10000000000000000000000011001000", b"00000000000000000000000000000000"),
	(b"00000000000001111110010111101011", b"00000000000001111110010100100011"), -- -2.8026e-43 + 7.25327e-40 = 7.25047e-40
	(b"01010110000010111011111011010011", b"00000000000000000000000000000000"),
	(b"10000000010011011100000000001101", b"01010110000010111011111011010011"), -- 3.84129e+13 + -7.14023e-39 = 3.84129e+13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100101111010010000001", b"11111111100000000000000000000000"), -- -inf + 1.74075e-39 = -inf
	(b"10101000001100110001000100101001", b"00000000000000000000000000000000"),
	(b"00000000010111001001000011111001", b"10101000001100110001000100101001"), -- -9.94022e-15 + 8.50087e-39 = -9.94022e-15
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110010000010001011110", b"11111111100000000000000000000000"), -- -inf + -8.17493e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000000011110111001101", b"11111111100000000000000000000000"), -- -inf + 2.96091e-39 = -inf
	(b"10011110000000010110000110101000", b"00000000000000000000000000000000"),
	(b"00000000001000101001011100000000", b"10011110000000010110000110101000"), -- -6.8494e-21 + 3.17658e-39 = -6.8494e-21
	(b"01010110000000111101001011111100", b"00000000000000000000000000000000"),
	(b"00000000010001000000001110100011", b"01010110000000111101001011111100"), -- 3.62355e+13 + 6.24612e-39 = 3.62355e+13
	(b"10100001011010000010111110010110", b"00000000000000000000000000000000"),
	(b"00000000001101011101100101101100", b"10100001011010000010111110010110"), -- -7.86676e-19 + 4.94528e-39 = -7.86676e-19
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100100101111110010100", b"00000000000100100101111110010100"), -- 0 + 1.68733e-39 = 1.68733e-39
	(b"10111010100010010101011010100111", b"00000000000000000000000000000000"),
	(b"10000000000100110011110110010001", b"10111010100010010101011010100111"), -- -0.00104781 + -1.76696e-39 = -0.00104781
	(b"00000010111100010100111010010110", b"00000000000000000000000000000000"),
	(b"00000000000010001010000001111010", b"00000010111100011101100010011110"), -- 3.54569e-37 + 7.92252e-40 = 3.55361e-37
	(b"10100110010100011001011110100001", b"00000000000000000000000000000000"),
	(b"00000000010010101010001110000100", b"10100110010100011001011110100001"), -- -7.27169e-16 + 6.85449e-39 = -7.27169e-16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110111001001000000001", b"10000000010110111001001000000001"), -- 0 + -8.40941e-39 = -8.40941e-39
	(b"10111011001101110110111110000111", b"00000000000000000000000000000000"),
	(b"00000000001010110111001001110000", b"10111011001101110110111110000111"), -- -0.00279901 + 3.98998e-39 = -0.00279901
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010111101011110110000", b"00000000001010111101011110110000"), -- 0 + 4.0263e-39 = 4.0263e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001011111101001011010101", b"00000000001011111101001011010101"), -- 0 + 4.3919e-39 = 4.3919e-39
	(b"00000001001101101001111000100110", b"00000000000000000000000000000000"),
	(b"10000000000011110000101101011101", b"00000001001011110001100001111000"), -- 3.35416e-38 + -1.38161e-39 = 3.216e-38
	(b"10100001111111111001100101011011", b"00000000000000000000000000000000"),
	(b"00000000011100011011010010100010", b"10100001111111111001100101011011"), -- -1.73201e-18 + 1.04422e-38 = -1.73201e-18
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010111000111011001010000", b"00000000010111000111011001010000"), -- -0 + 8.49131e-39 = 8.49131e-39
	(b"01101101011010000010000101010010", b"00000000000000000000000000000000"),
	(b"00000000010010100011011011000100", b"01101101011010000010000101010010"), -- 4.49005e+27 + 6.81547e-39 = 4.49005e+27
	(b"01101100001010111000010101001101", b"00000000000000000000000000000000"),
	(b"10000000010011001111010011000010", b"01101100001010111000010101001101"), -- 8.29423e+26 + -7.0673e-39 = 8.29423e+26
	(b"00111000111011110100000000001110", b"00000000000000000000000000000000"),
	(b"00000000010111101111000101010010", b"00111000111011110100000000001110"), -- 0.000114083 + 8.71911e-39 = 0.000114083
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001011101011010100110100", b"01111111100000000000000000000000"), -- inf + -4.28944e-39 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000101000111110000011011", b"11111111100000000000000000000000"), -- -inf + -1.88123e-39 = -inf
	(b"10100001000100111111110101001010", b"00000000000000000000000000000000"),
	(b"00000000010100000111100110011011", b"10100001000100111111110101001010"), -- -5.01408e-19 + 7.39046e-39 = -5.01408e-19
	(b"11110100010001010111110111001111", b"00000000000000000000000000000000"),
	(b"00000000010110001111000011001111", b"11110100010001010111110111001111"), -- -6.25875e+31 + 8.16791e-39 = -6.25875e+31
	(b"10000101010111110000011001000110", b"00000000000000000000000000000000"),
	(b"00000000000101101100010010101111", b"10000101010111101111101011100100"), -- -1.04866e-35 + 2.09094e-39 = -1.04845e-35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001011000011110011111001", b"11111111100000000000000000000000"), -- -inf + -4.06263e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100000011110011001000", b"01111111100000000000000000000000"), -- inf + -1.03074e-38 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001100011110000100010100", b"10000000001100011110000100010100"), -- 0 + -4.58068e-39 = -4.58068e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110100110011111100001", b"01111111100000000000000000000000"), -- inf + -8.30246e-39 = inf
	(b"10101101011111100000001010111100", b"00000000000000000000000000000000"),
	(b"00000000010111011001000010001010", b"10101101011111100000001010111100"), -- -1.44388e-11 + 8.59255e-39 = -1.44388e-11
	(b"10011010111110001000000111110110", b"00000000000000000000000000000000"),
	(b"00000000010110010010011011001101", b"10011010111110001000000111110110"), -- -1.0278e-22 + 8.18728e-39 = -1.0278e-22
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011000100011010010011", b"11111111100000000000000000000000"), -- -inf + -1.12734e-39 = -inf
	(b"01010101010011100000110000111001", b"00000000000000000000000000000000"),
	(b"00000000011111010100101001001010", b"01010101010011100000110000111001"), -- 1.41595e+13 + 1.15061e-38 = 1.41595e+13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010110111100000001000000", b"11111111100000000000000000000000"), -- -inf + 8.426e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000100000100000000010", b"01111111100000000000000000000000"), -- inf + -1.86544e-40 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000111001000100111011111", b"01111111100000000000000000000000"), -- inf + -2.62085e-39 = inf
	(b"10010101110111111010101010100110", b"00000000000000000000000000000000"),
	(b"10000000011110100000010001010110", b"10010101110111111010101010100110"), -- -9.03382e-26 + -1.12055e-38 = -9.03382e-26
	(b"01011101111111110001010011110110", b"00000000000000000000000000000000"),
	(b"00000000011111110101100011101110", b"01011101111111110001010011110110"), -- 2.29757e+18 + 1.1695e-38 = 2.29757e+18
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011010110010110111000101", b"10000000011010110010110111000101"), -- -0 + -9.84282e-39 = -9.84282e-39
	(b"10011101101110011111001000110000", b"00000000000000000000000000000000"),
	(b"10000000010001010100111111000011", b"10011101101110011111001000110000"), -- -4.92195e-21 + -6.36526e-39 = -4.92195e-21
	(b"10100000011101101101101101100000", b"00000000000000000000000000000000"),
	(b"10000000001000011101101011011010", b"10100000011101101101101101100000"), -- -2.09096e-19 + -3.10908e-39 = -2.09096e-19
	(b"10000110000100100011111011110010", b"00000000000000000000000000000000"),
	(b"10000000000100000110001111000110", b"10000110000100100100000011111110"), -- -2.75058e-35 + -1.50516e-39 = -2.75073e-35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000111110010100100101010", b"11111111100000000000000000000000"), -- -inf + -2.86167e-39 = -inf
	(b"00001100001101110111000101100001", b"00000000000000000000000000000000"),
	(b"00000000010100010011110011101111", b"00001100001101110111000101100010"), -- 1.41319e-31 + 7.46053e-39 = 1.41319e-31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001111000110110100101", b"00000000011001111000110110100101"), -- -0 + 9.50987e-39 = 9.50987e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001110010010101001011", b"00000000000001110010010101001011"), -- -0 + 6.56227e-40 = 6.56227e-40
	(b"10101110010110110010111000010111", b"00000000000000000000000000000000"),
	(b"00000000001100111101101011000011", b"10101110010110110010111000010111"), -- -4.98358e-11 + 4.76209e-39 = -4.98358e-11
	(b"11011010000101000110110000110011", b"00000000000000000000000000000000"),
	(b"00000000010101111100101101100101", b"11011010000101000110110000110011"), -- -1.04443e+16 + 8.06265e-39 = -1.04443e+16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000001110100010111111", b"00000000001000001110100010111111"), -- 0 + 3.02223e-39 = 3.02223e-39
	(b"10000111100101011010110011111001", b"00000000000000000000000000000000"),
	(b"00000000010010110001000100111011", b"10000111100101011010101111001101"), -- -2.25207e-34 + 6.89384e-39 = -2.252e-34
	(b"00101011010111000110011110111011", b"00000000000000000000000000000000"),
	(b"10000000000000100111110111110001", b"00101011010111000110011110111011"), -- 7.83037e-13 + -2.2885e-40 = 7.83037e-13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000001000101111011110111", b"11111111100000000000000000000000"), -- -inf + -4.01409e-40 = -inf
	(b"11010110010011011101010000010000", b"00000000000000000000000000000000"),
	(b"10000000010010001110011000100111", b"11010110010011011101010000010000"), -- -5.65777e+13 + -6.69472e-39 = -5.65777e+13
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011001101010011011100010", b"00000000011001101010011011100010"), -- 0 + 9.42709e-39 = 9.42709e-39
	(b"00000000000000000000000000000011", b"00000000000000000000000000000000"),
	(b"10000000000010000101000110101011", b"10000000000010000101000110101000"), -- 4.2039e-45 + -7.63981e-40 = -7.63977e-40
	(b"00101100011101111010001100101110", b"00000000000000000000000000000000"),
	(b"00000000000010000111110011011011", b"00101100011101111010001100101110"), -- 3.51914e-12 + 7.79474e-40 = 3.51914e-12
	(b"10000000000000000000000110101011", b"00000000000000000000000000000000"),
	(b"10000000011111010111101010001101", b"10000000011111010111110000111000"), -- -5.98354e-43 + -1.15234e-38 = -1.1524e-38
	(b"10111011010100110110001111000101", b"00000000000000000000000000000000"),
	(b"00000000000110100101100110011101", b"10111011010100110110001111000101"), -- -0.00322555 + 2.41987e-39 = -0.00322555
	(b"01000010100010010100001011011100", b"00000000000000000000000000000000"),
	(b"00000000001110001011010010110111", b"01000010100010010100001011011100"), -- 68.6306 + 5.20762e-39 = 68.6306
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001111000111110100100011", b"00000000001111000111110100100011"), -- 0 + 5.55502e-39 = 5.55502e-39
	(b"11110010000001011011001000000111", b"00000000000000000000000000000000"),
	(b"10000000010000000010110101010010", b"11110010000001011011001000000111"), -- -2.64811e+30 + -5.89373e-39 = -2.64811e+30
	(b"01101000001111001101111000000010", b"00000000000000000000000000000000"),
	(b"00000000001111111101000100001101", b"01101000001111001101111000000010"), -- 3.5676e+24 + 5.86063e-39 = 3.5676e+24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101010111011000011011", b"10000000001101010111011000011011"), -- -0 + -4.90965e-39 = -4.90965e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000011000011011010001", b"10000000011000011000011011010001"), -- -0 + -8.95641e-39 = -8.95641e-39
	(b"00001111000111111010011011010000", b"00000000000000000000000000000000"),
	(b"00000000010110001110111000101101", b"00001111000111111010011011010000"), -- 7.87143e-30 + 8.16697e-39 = 7.87143e-30
	(b"01101001010110000000000101100010", b"00000000000000000000000000000000"),
	(b"10000000010000100010011100101010", b"01101001010110000000000101100010"), -- 1.63209e+25 + -6.07519e-39 = 1.63209e+25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101110011010001010111", b"11111111100000000000000000000000"), -- -inf + -5.06973e-39 = -inf
	(b"10000011111110111011100011100101", b"00000000000000000000000000000000"),
	(b"00000000010011000101000101100100", b"10000011111110101000011110011111"), -- -1.47949e-36 + 7.0087e-39 = -1.47248e-36
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110001101110000110100", b"01111111100000000000000000000000"), -- inf + -1.10993e-38 = inf
	(b"01101111110100010011000011110111", b"00000000000000000000000000000000"),
	(b"00000000011010100111110101110111", b"01101111110100010011000011110111"), -- 1.29483e+29 + 9.77957e-39 = 1.29483e+29
	(b"10011001101101101011010111111110", b"00000000000000000000000000000000"),
	(b"10000000000110110001010101110100", b"10011001101101101011010111111110"), -- -1.88919e-23 + -2.48725e-39 = -1.88919e-23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001011110001101010111001", b"10000000001011110001101010111001"), -- 0 + -4.32585e-39 = -4.32585e-39
	(b"00111011001100101000010111111100", b"00000000000000000000000000000000"),
	(b"00000000011010101000001100100110", b"00111011001100101000010111111100"), -- 0.00272405 + 9.78161e-39 = 0.00272405
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101111010000000001000", b"01111111100000000000000000000000"), -- inf + -5.10836e-39 = inf
	(b"11111000110110001101101010111110", b"00000000000000000000000000000000"),
	(b"00000000000011101001111111100101", b"11111000110110001101101010111110"), -- -3.51866e+34 + 1.34306e-39 = -3.51866e+34
	(b"00000000000000000000001101001000", b"00000000000000000000000000000000"),
	(b"10000000011001001000011101110011", b"10000000011001001000010000101011"), -- 1.17709e-42 + -9.23214e-39 = -9.23096e-39
	(b"01100000111000000011001100010010", b"00000000000000000000000000000000"),
	(b"10000000000111000100101001111110", b"01100000111000000011001100010010"), -- 1.29242e+20 + -2.59812e-39 = 1.29242e+20
	(b"01111000000110100110111011000001", b"00000000000000000000000000000000"),
	(b"00000000010111100001000111010000", b"01111000000110100110111011000001"), -- 1.25291e+34 + 8.63893e-39 = 1.25291e+34
	(b"10111111001110111110101101010000", b"00000000000000000000000000000000"),
	(b"00000000011011011111101010100010", b"10111111001110111110101101010000"), -- -0.734059 + 1.01e-38 = -0.734059
	(b"10101000001011011010111110101100", b"00000000000000000000000000000000"),
	(b"00000000011001110011110100110011", b"10101000001011011010111110101100"), -- -9.64152e-15 + 9.48101e-39 = -9.64152e-15
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101100001100001100011", b"11111111100000000000000000000000"), -- -inf + 1.08453e-38 = -inf
	(b"11110010100010010010010001000101", b"00000000000000000000000000000000"),
	(b"10000000011110000101010000111000", b"11110010100010010010010001000101"), -- -5.43274e+30 + -1.10505e-38 = -5.43274e+30
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001100001001000001111100", b"01111111100000000000000000000000"), -- inf + 4.45994e-39 = inf
	(b"00100011100000011110010111010000", b"00000000000000000000000000000000"),
	(b"00000000011001011011000000010111", b"00100011100000011110010111010000"), -- 1.40835e-17 + 9.33855e-39 = 1.40835e-17
	(b"10110000000100000011010001011001", b"00000000000000000000000000000000"),
	(b"10000000010011101111100010010111", b"10110000000100000011010001011001"), -- -5.24613e-10 + -7.25235e-39 = -5.24613e-10
	(b"10010010111101000000000001100101", b"00000000000000000000000000000000"),
	(b"00000000010110001000011111110001", b"10010010111101000000000001100101"), -- -1.53987e-27 + 8.13029e-39 = -1.53987e-27
	(b"11000110100111101100101110011001", b"00000000000000000000000000000000"),
	(b"10000000010100101110000110000100", b"11000110100111101100101110011001"), -- -20325.8 + -7.61141e-39 = -20325.8
	(b"10100111100111001011000101110000", b"00000000000000000000000000000000"),
	(b"00000000011101101100111001101011", b"10100111100111001011000101110000"), -- -4.34911e-15 + 1.09106e-38 = -4.34911e-15
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010010011110000010010", b"10000000000010010011110000010010"), -- 0 + -8.48069e-40 = -8.48069e-40
	(b"11101100010101001011000111111111", b"00000000000000000000000000000000"),
	(b"10000000010100101011010111010001", b"11101100010101001011000111111111"), -- -1.02853e+27 + -7.59573e-39 = -1.02853e+27
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001101001101001011111001", b"01111111100000000000000000000000"), -- inf + -4.85113e-39 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001000111000000010111011", b"01111111100000000000000000000000"), -- inf + 3.26042e-39 = inf
	(b"01011010000111001100001000100110", b"00000000000000000000000000000000"),
	(b"00000000011001110010100001110001", b"01011010000111001100001000100110"), -- 1.10309e+16 + 9.47356e-39 = 1.10309e+16
	(b"01100000001111001001001100101110", b"00000000000000000000000000000000"),
	(b"00000000011101110101100111111000", b"01100000001111001001001100101110"), -- 5.4353e+19 + 1.09607e-38 = 5.4353e+19
	(b"11111010000101100100111101001110", b"00000000000000000000000000000000"),
	(b"00000000011010000100011101111101", b"11111010000101100100111101001110"), -- -1.95113e+35 + 9.57654e-39 = -1.95113e+35
	(b"10011011011101001101010101110101", b"00000000000000000000000000000000"),
	(b"00000000011011010000100001110000", b"10011011011101001101010101110101"), -- -2.02522e-22 + 1.00131e-38 = -2.02522e-22
	(b"11111001010000000101100001010101", b"00000000000000000000000000000000"),
	(b"10000000000111011101100011100101", b"11111001010000000101100001010101"), -- -6.24195e+34 + -2.74104e-39 = -6.24195e+34
	(b"10111111101111001111011001010111", b"00000000000000000000000000000000"),
	(b"00000000000111111100011001010110", b"10111111101111001111011001010111"), -- -1.47627 + 2.91805e-39 = -1.47627
	(b"01000001110101100101100000000101", b"00000000000000000000000000000000"),
	(b"00000000010001000110000111100010", b"01000001110101100101100000000101"), -- 26.793 + 6.27993e-39 = 26.793
	(b"00000000000000000000000000111001", b"00000000000000000000000000000000"),
	(b"00000000011011110000101011101101", b"00000000011011110000101100100110"), -- 7.9874e-44 + 1.01977e-38 = 1.01977e-38
	(b"10000010101010101111011101010100", b"00000000000000000000000000000000"),
	(b"10000000011010010010010010100000", b"10000010101100011000100110011110"), -- -2.51212e-37 + -9.65587e-39 = -2.60868e-37
	(b"11001000100011101101101011010100", b"00000000000000000000000000000000"),
	(b"10000000001101110010000001111101", b"11001000100011101101101011010100"), -- -292567 + -5.06261e-39 = -292567
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010001100100001011100", b"10000000001010001100100001011100"), -- -0 + -3.7453e-39 = -3.7453e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011111101101001011011001", b"11111111100000000000000000000000"), -- -inf + -1.16469e-38 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101111100001001101011", b"00000000011101111100001001101011"), -- 0 + 1.09982e-38 = 1.09982e-38
	(b"01000000011101001110010010110010", b"00000000000000000000000000000000"),
	(b"10000000011000010111110110101110", b"01000000011101001110010010110010"), -- 3.82646 + -8.95313e-39 = 3.82646
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001101101010000000110101", b"01111111100000000000000000000000"), -- inf + 5.01659e-39 = inf
	(b"10111101110001000100111101101110", b"00000000000000000000000000000000"),
	(b"00000000000011000000001000000001", b"10111101110001000100111101101110"), -- -0.0958546 + 1.10274e-39 = -0.0958546
	(b"01111101100000000101000011001011", b"00000000000000000000000000000000"),
	(b"10000000001111110010110101000000", b"01111101100000000101000011001011"), -- 2.13201e+37 + -5.80187e-39 = 2.13201e+37
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010010110101000100000101", b"00000000010010110101000100000101"), -- 0 + 6.91673e-39 = 6.91673e-39
	(b"11101110100011011011100101111111", b"00000000000000000000000000000000"),
	(b"00000000011001111011000000110101", b"11101110100011011011100101111111"), -- -2.19308e+28 + 9.52227e-39 = -2.19308e+28
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010101110010010100110111", b"00000000010101110010010100110111"), -- -0 + 8.00304e-39 = 8.00304e-39
	(b"10100010101011010111000011111010", b"00000000000000000000000000000000"),
	(b"10000000000011111110011110011101", b"10100010101011010111000011111010"), -- -4.70114e-18 + -1.46062e-39 = -4.70114e-18
	(b"00111111110010011101110010011100", b"00000000000000000000000000000000"),
	(b"00000000010011000111111011110100", b"00111111110010011101110010011100"), -- 1.57704 + 7.02504e-39 = 1.57704
	(b"00111011101100100000010001101010", b"00000000000000000000000000000000"),
	(b"00000000011111111010001000000010", b"00111011101100100000010001101010"), -- 0.00543266 + 1.17212e-38 = 0.00543266
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010111011101000010000111", b"10000000010111011101000010000111"), -- -0 + -8.61551e-39 = -8.61551e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110111011011101101010", b"01111111100000000000000000000000"), -- inf + -1.13616e-38 = inf
	(b"10111101111011110000111010011110", b"00000000000000000000000000000000"),
	(b"10000000010001111100000010100000", b"10111101111011110000111010011110"), -- -0.116727 + -6.58942e-39 = -0.116727
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010101100101001101101011", b"11111111100000000000000000000000"), -- -inf + 7.92778e-39 = -inf
	(b"11110010010101100010011011110111", b"00000000000000000000000000000000"),
	(b"10000000011111010111010011110111", b"11110010010101100010011011110111"), -- -4.24172e+30 + -1.15214e-38 = -4.24172e+30
	(b"00011001100111111011001010101111", b"00000000000000000000000000000000"),
	(b"10000000001010100100110110000011", b"00011001100111111011001010101111"), -- 1.65124e-23 + -3.8849e-39 = 1.65124e-23
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011101000101110100001110", b"11111111100000000000000000000000"), -- -inf + 1.06863e-38 = -inf
	(b"11101100100100001000000101011000", b"00000000000000000000000000000000"),
	(b"00000000011000001100000111110001", b"11101100100100001000000101011000"), -- -1.39757e+27 + 8.88578e-39 = -1.39757e+27
	(b"10011011010010010100001011011100", b"00000000000000000000000000000000"),
	(b"10000000000001111110000010000011", b"10011011010010010100001011011100"), -- -1.66479e-22 + -7.23388e-40 = -1.66479e-22
	(b"00000000000000000000000001101011", b"00000000000000000000000000000000"),
	(b"00000000001110000101101101111000", b"00000000001110000101101111100011"), -- 1.49939e-43 + 5.1756e-39 = 5.17575e-39
	(b"11010011001100000010000011011110", b"00000000000000000000000000000000"),
	(b"10000000011001111011100001111101", b"11010011001100000010000011011110"), -- -7.56466e+11 + -9.52524e-39 = -7.56466e+11
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000100001101000000000110", b"00000000000100001101000000000110"), -- -0 + 1.54399e-39 = 1.54399e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001001100001001110011", b"01111111100000000000000000000000"), -- inf + 6.31457e-39 = inf
	(b"00000000000000010010001111100000", b"00000000000000000000000000000000"),
	(b"10000000010011001001011100000100", b"10000000010010110111001100100100"), -- 1.04705e-40 + -7.03367e-39 = -6.92897e-39
	(b"01001001101100110010011011001011", b"00000000000000000000000000000000"),
	(b"00000000000000100101100110110111", b"01001001101100110010011011001011"), -- 1.46761e+06 + 2.15855e-40 = 1.46761e+06
	(b"01001011000110101101101100010001", b"00000000000000000000000000000000"),
	(b"10000000000000010010000001000011", b"01001011000110101101101100010001"), -- 1.01486e+07 + -1.03409e-40 = 1.01486e+07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000110000001110100010100", b"11111111100000000000000000000000"), -- -inf + -2.21448e-39 = -inf
	(b"10110010000110101000100101110010", b"00000000000000000000000000000000"),
	(b"10000000001100011011110001000000", b"10110010000110101000100101110010"), -- -8.99523e-09 + -4.56747e-39 = -8.99523e-09
	(b"00000101101111001110100010101010", b"00000000000000000000000000000000"),
	(b"00000000010000100100111000110110", b"00000101101111001111100100111110"), -- 1.77649e-35 + 6.0892e-39 = 1.7771e-35
	(b"00011010110011100011001101110000", b"00000000000000000000000000000000"),
	(b"10000000011101101011011011111100", b"00011010110011100011001101110000"), -- 8.52827e-23 + -1.09022e-38 = 8.52827e-23
	(b"01011010010100000100010111110110", b"00000000000000000000000000000000"),
	(b"00000000011111010011101100110000", b"01011010010100000100010111110110"), -- 1.46559e+16 + 1.15007e-38 = 1.46559e+16
	(b"10110000100101011111110000101100", b"00000000000000000000000000000000"),
	(b"00000000001001010011100101000010", b"10110000100101011111110000101100"), -- -1.09128e-09 + 3.41845e-39 = -1.09128e-09
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001100011110010010011", b"11111111100000000000000000000000"), -- -inf + -3.51148e-39 = -inf
	(b"01010010100110000101011111110000", b"00000000000000000000000000000000"),
	(b"00000000000111111100110101111100", b"01010010100110000101011111110000"), -- 3.27155e+11 + 2.92061e-39 = 3.27155e+11
	(b"00101110000010101101100100010000", b"00000000000000000000000000000000"),
	(b"10000000001010111110010011001011", b"00101110000010101101100100010000"), -- 3.15704e-11 + -4.031e-39 = 3.15704e-11
	(b"01101111110010001010011000000001", b"00000000000000000000000000000000"),
	(b"10000000000010000011100010101010", b"01101111110010001010011000000001"), -- 1.24195e+29 + -7.55011e-40 = 1.24195e+29
	(b"00010011111111001000000001010011", b"00000000000000000000000000000000"),
	(b"10000000010101111010011000011011", b"00010011111111001000000001010011"), -- 6.37403e-27 + -8.04928e-39 = 6.37403e-27
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000010110010111110100", b"10000000000000010110010111110100"), -- 0 + -1.28409e-40 = -1.28409e-40
	(b"10010111101100010000000110001110", b"00000000000000000000000000000000"),
	(b"00000000010011111110001101101000", b"10010111101100010000000110001110"), -- -1.14387e-24 + 7.33658e-39 = -1.14387e-24
	(b"00000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"10000000000111110101010111010010", b"10000000000111110101010111010001"), -- 1.4013e-45 + -2.87769e-39 = -2.87769e-39
	(b"10101100000001011010101010100101", b"00000000000000000000000000000000"),
	(b"00000000010110101100111010101100", b"10101100000001011010101010100101"), -- -1.89952e-12 + 8.33933e-39 = -1.89952e-12
	(b"01010111100000101100100001000010", b"00000000000000000000000000000000"),
	(b"10000000000001011110011101000011", b"01010111100000101100100001000010"), -- 2.87593e+14 + -5.42139e-40 = 2.87593e+14
	(b"11010000110000010100110110101010", b"00000000000000000000000000000000"),
	(b"10000000011001101010001010010111", b"11010000110000010100110110101010"), -- -2.59447e+10 + -9.42555e-39 = -2.59447e+10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000111001000110110101110", b"11111111100000000000000000000000"), -- -inf + 2.62222e-39 = -inf
	(b"10011100011011001110101001111110", b"00000000000000000000000000000000"),
	(b"10000000000101101011001000100000", b"10011100011011001110101001111110"), -- -7.83889e-22 + -2.08428e-39 = -7.83889e-22
	(b"00010111010001000101000010011111", b"00000000000000000000000000000000"),
	(b"00000000000110011001101101010011", b"00010111010001000101000010011111"), -- 6.34328e-25 + 2.35161e-39 = 6.34328e-25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001011100100110111011111", b"11111111100000000000000000000000"), -- -inf + -4.25237e-39 = -inf
	(b"01010001101111000011110110110001", b"00000000000000000000000000000000"),
	(b"10000000000110001000100110100010", b"01010001101111000011110110110001"), -- 1.01061e+11 + -2.25343e-39 = 1.01061e+11
	(b"10100010111100110100001101111101", b"00000000000000000000000000000000"),
	(b"10000000011111001101010111010110", b"10100010111100110100001101111101"), -- -6.59367e-18 + -1.14643e-38 = -6.59367e-18
	(b"01110101110110100111011110010101", b"00000000000000000000000000000000"),
	(b"10000000011100001100010010100011", b"01110101110110100111011110010101"), -- 5.5388e+32 + -1.03561e-38 = 5.5388e+32
	(b"10001011110111111110000001001100", b"00000000000000000000000000000000"),
	(b"00000000000100101101111101110111", b"10001011110111111110000001001100"), -- -8.6234e-32 + 1.7332e-39 = -8.6234e-32
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011000101001000101011111", b"01111111100000000000000000000000"), -- inf + -9.05203e-39 = inf
	(b"01101110010100100001010110101011", b"00000000000000000000000000000000"),
	(b"00000000011111001111110001011001", b"01101110010100100001010110101011"), -- 1.62545e+28 + 1.14781e-38 = 1.62545e+28
	(b"10110010011011101011110001100100", b"00000000000000000000000000000000"),
	(b"10000000011010010001001101001110", b"10110010011011101011110001100100"), -- -1.38963e-08 + -9.64965e-39 = -1.38963e-08
	(b"00000100110100111100100011101110", b"00000000000000000000000000000000"),
	(b"10000000001000000101010011000001", b"00000100110100111010100010011001"), -- 4.97904e-36 + -2.96914e-39 = 4.97607e-36
	(b"10001111010001110010011111010011", b"00000000000000000000000000000000"),
	(b"10000000011110001110010001110110", b"10001111010001110010011111010011"), -- -9.81913e-30 + -1.11022e-38 = -9.81913e-30
	(b"10101000101001011011101000000100", b"00000000000000000000000000000000"),
	(b"10000000000101000100111100001101", b"10101000101001011011101000000100"), -- -1.83994e-14 + -1.86507e-39 = -1.83994e-14
	(b"01101001001011011010111001011110", b"00000000000000000000000000000000"),
	(b"00000000011010100100110101001011", b"01101001001011011010111001011110"), -- 1.3123e+25 + 9.76229e-39 = 1.3123e+25
	(b"10110010111011011101011011011100", b"00000000000000000000000000000000"),
	(b"10000000010100110101111111111000", b"10110010111011011101011011011100"), -- -2.76881e-08 + -7.65677e-39 = -2.76881e-08
	(b"01001001111001001010001101100001", b"00000000000000000000000000000000"),
	(b"00000000010111010011110110011010", b"01001001111001001010001101100001"), -- 1.873e+06 + 8.5628e-39 = 1.873e+06
	(b"01010000111100100011100010110010", b"00000000000000000000000000000000"),
	(b"10000000001011110011000111101101", b"01010000111100100011100010110010"), -- 3.25104e+10 + -4.33418e-39 = 3.25104e+10
	(b"01001100110011100110011100000110", b"00000000000000000000000000000000"),
	(b"00000000001111000010111001110011", b"01001100110011100110011100000110"), -- 1.08214e+08 + 5.52679e-39 = 1.08214e+08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010110011100001000111", b"01111111100000000000000000000000"), -- inf + -1.03038e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010111111001101010101101", b"00000000010111111001101010101101"), -- 0 + 8.77986e-39 = 8.77986e-39
	(b"10101000111100001010011001110100", b"00000000000000000000000000000000"),
	(b"10000000011111111100101001111111", b"10101000111100001010011001110100"), -- -2.67175e-14 + -1.17357e-38 = -2.67175e-14
	(b"11011010100101110111011110010001", b"00000000000000000000000000000000"),
	(b"00000000011111011001101100001101", b"11011010100101110111011110010001"), -- -2.13171e+16 + 1.15351e-38 = -2.13171e+16
	(b"10011000010011000111111000001101", b"00000000000000000000000000000000"),
	(b"00000000001000000010111100011000", b"10011000010011000111111000001101"), -- -2.643e-24 + 2.95563e-39 = -2.643e-24
	(b"00000000000000000001010111010101", b"00000000000000000000000000000000"),
	(b"10000000011000000000011111100100", b"10000000010111111111001000001111"), -- 7.83186e-42 + -8.81904e-39 = -8.81121e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010110010111001111010010", b"11111111100000000000000000000000"), -- -inf + -8.21491e-39 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010101100101101101111100", b"10000000010101100101101101111100"), -- 0 + -7.93067e-39 = -7.93067e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011010110111111001110100", b"10000000011010110111111001110100"), -- -0 + -9.87176e-39 = -9.87176e-39
	(b"10101110100001010000110100010100", b"00000000000000000000000000000000"),
	(b"00000000011000101011101110000011", b"10101110100001010000110100010100"), -- -6.05046e-11 + 9.06715e-39 = -6.05046e-11
	(b"00111110001100100000011001000101", b"00000000000000000000000000000000"),
	(b"10000000001110100001010000011001", b"00111110001100100000011001000101"), -- 0.173852 + -5.33367e-39 = 0.173852
	(b"00010010101100100111111000000000", b"00000000000000000000000000000000"),
	(b"00000000001010111001111111101000", b"00010010101100100111111000000000"), -- 1.12644e-27 + 4.00629e-39 = 1.12644e-27
	(b"11010001000000111110111011000101", b"00000000000000000000000000000000"),
	(b"00000000010011011000111100101000", b"11010001000000111110111011000101"), -- -3.54154e+10 + 7.12269e-39 = -3.54154e+10
	(b"10110011110110011110010110000010", b"00000000000000000000000000000000"),
	(b"00000000010100000001110101011000", b"10110011110110011110010110000010"), -- -1.01466e-07 + 7.35737e-39 = -1.01466e-07
	(b"01010101101110111000111100110000", b"00000000000000000000000000000000"),
	(b"00000000001110001101111001100011", b"01010101101110111000111100110000"), -- 2.5778e+13 + 5.22257e-39 = 2.5778e+13
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011100110111100111010", b"10000000000011100110111100111010"), -- 0 + -1.3256e-39 = -1.3256e-39
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"10000000001100011000000000111111", b"10000000001100011000000001000000"), -- -1.4013e-45 + -4.54595e-39 = -4.54595e-39
	(b"11100110000110011110001010000100", b"00000000000000000000000000000000"),
	(b"00000000000001000111000110000111", b"11100110000110011110001010000100"), -- -1.81675e+23 + 4.08068e-40 = -1.81675e+23
	(b"10100111100110000111010101011101", b"00000000000000000000000000000000"),
	(b"10000000010111000111010100110110", b"10100111100110000111010101011101"), -- -4.23157e-15 + -8.49091e-39 = -4.23157e-15
	(b"11100001110111101110010001110110", b"00000000000000000000000000000000"),
	(b"00000000001111100100110100110011", b"11100001110111101110010001110110"), -- -5.13955e+20 + 5.72149e-39 = -5.13955e+20
	(b"10001111101001011100001100001001", b"00000000000000000000000000000000"),
	(b"00000000000011111111000100001001", b"10001111101001011100001100001001"), -- -1.63454e-29 + 1.464e-39 = -1.63454e-29
	(b"10101101111001001111101000101111", b"00000000000000000000000000000000"),
	(b"10000000010001001011001000101011", b"10101101111001001111101000101111"), -- -2.60317e-11 + -6.30873e-39 = -2.60317e-11
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011100110001010101101101", b"01111111100000000000000000000000"), -- inf + 1.05688e-38 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110010111000110010101", b"10000000001110010111000110010101"), -- -0 + -5.27537e-39 = -5.27537e-39
	(b"01010001000001111000010110110011", b"00000000000000000000000000000000"),
	(b"10000000000100001010100010010101", b"01010001000001111000010110110011"), -- 3.6379e+10 + -1.52984e-39 = 3.6379e+10
	(b"11111101111100111000011010111000", b"00000000000000000000000000000000"),
	(b"00000000000000110000010100001111", b"11111101111100111000011010111000"), -- -4.04627e+37 + 2.77321e-40 = -4.04627e+37
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001010101100111011110", b"00000000000001010101100111011110"), -- 0 + 4.91416e-40 = 4.91416e-40
	(b"11101111001000101100011001000010", b"00000000000000000000000000000000"),
	(b"00000000011110111110011010100000", b"11101111001000101100011001000010"), -- -5.03763e+28 + 1.13785e-38 = -5.03763e+28
	(b"01011000010111100001011001001011", b"00000000000000000000000000000000"),
	(b"10000000011100110001010010001011", b"01011000010111100001011001001011"), -- 9.76749e+14 + -1.05685e-38 = 9.76749e+14
	(b"01010110100000101001100000101101", b"00000000000000000000000000000000"),
	(b"10000000001010010000100011111100", b"01010110100000101001100000101101"), -- 7.17951e+13 + -3.76848e-39 = 7.17951e+13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000010011100110010101101", b"01111111100000000000000000000000"), -- inf + -8.99943e-40 = inf
	(b"00101110000001101101011001001000", b"00000000000000000000000000000000"),
	(b"00000000000100001001011110100101", b"00101110000001101101011001001000"), -- 3.06584e-11 + 1.52377e-39 = 3.06584e-11
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000010001110001010001001000", b"01111111100000000000000000000000"), -- inf + -6.5276e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001001001110011101101100", b"10000000001001001110011101101100"), -- 0 + -3.3891e-39 = -3.3891e-39
	(b"10111110000000000110011001110001", b"00000000000000000000000000000000"),
	(b"10000000000101000101111110101010", b"10111110000000000110011001110001"), -- -0.125391 + -1.87103e-39 = -0.125391
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001010010101101011110011", b"10000000001010010101101011110011"), -- -0 + -3.79788e-39 = -3.79788e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001110110011011101000111", b"10000000001110110011011101000111"), -- -0 + -5.43812e-39 = -5.43812e-39
	(b"10011110101010001111101100010100", b"00000000000000000000000000000000"),
	(b"00000000010000100011101000010001", b"10011110101010001111101100010100"), -- -1.78915e-20 + 6.08197e-39 = -1.78915e-20
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110010101111110011010", b"11111111100000000000000000000000"), -- -inf + 5.26892e-39 = -inf
	(b"10111011001001000011100010100111", b"00000000000000000000000000000000"),
	(b"10000000001100001111001111000101", b"10111011001001000011100010100111"), -- -0.00250582 + -4.49555e-39 = -0.00250582
	(b"10011001011001001100111010010000", b"00000000000000000000000000000000"),
	(b"10000000001000011010110010010000", b"10011001011001001100111010010000"), -- -1.1829e-23 + -3.09248e-39 = -1.1829e-23
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000011100101000011010100", b"01111111100000000000000000000000"), -- inf + -1.31469e-39 = inf
	(b"11111001011011101101001010011110", b"00000000000000000000000000000000"),
	(b"10000000011001000010111101111011", b"11111001011011101101001010011110"), -- -7.75024e+34 + -9.20058e-39 = -7.75024e+34
	(b"11110100010100111110110000110011", b"00000000000000000000000000000000"),
	(b"00000000001011101010111010000010", b"11110100010100111110110000110011"), -- -6.7161e+31 + 4.28703e-39 = -6.7161e+31
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000010000111111110110", b"01111111100000000000000000000000"), -- inf + 9.75612e-41 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000001010100100001011101", b"10000000000001010100100001011101"), -- 0 + -4.85137e-40 = -4.85137e-40
	(b"00110100011011001110111001011111", b"00000000000000000000000000000000"),
	(b"10000000001100000100111011111010", b"00110100011011001110111001011111"), -- 2.20659e-07 + -4.43644e-39 = 2.20659e-07
	(b"10100001110000000100100010101001", b"00000000000000000000000000000000"),
	(b"10000000000111111111101111101100", b"10100001110000000100100010101001"), -- -1.30297e-18 + -2.93727e-39 = -1.30297e-18
	(b"11100001001101001110011011011100", b"00000000000000000000000000000000"),
	(b"10000000000100111101100111110111", b"11100001001101001110011011011100"), -- -2.08566e+20 + -1.82307e-39 = -2.08566e+20
	(b"01110000101010001001110110110101", b"00000000000000000000000000000000"),
	(b"10000000000100111111110011101001", b"01110000101010001001110110110101"), -- 4.17473e+29 + -1.8356e-39 = 4.17473e+29
	(b"11000110100010100001111110001001", b"00000000000000000000000000000000"),
	(b"10000000000010111010000011010110", b"11000110100010100001111110001001"), -- -17679.8 + -1.06789e-39 = -17679.8
	(b"01000110111010110111101001001000", b"00000000000000000000000000000000"),
	(b"10000000011001101101100001110110", b"01000110111010110111101001001000"), -- 30141.1 + -9.44487e-39 = 30141.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001010110000010000010011", b"00000000001010110000010000010011"), -- 0 + 3.95039e-39 = 3.95039e-39
	(b"10010101101010110011110101111000", b"00000000000000000000000000000000"),
	(b"10000000001001001100011001000100", b"10010101101010110011110101111000"), -- -6.91633e-26 + -3.3772e-39 = -6.91633e-26
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011100011001011101000000", b"00000000011100011001011101000000"), -- 0 + 1.04317e-38 = 1.04317e-38
	(b"00111100000100001011010000000000", b"00000000000000000000000000000000"),
	(b"10000000011001110010101010111101", b"00111100000100001011010000000000"), -- 0.00883198 + -9.47439e-39 = 0.00883198
	(b"10101110000001011100101111000000", b"00000000000000000000000000000000"),
	(b"00000000000110111000101100001010", b"10101110000001011100101111000000"), -- -3.04217e-11 + 2.52944e-39 = -3.04217e-11
	(b"10010111111111001111000001011110", b"00000000000000000000000000000000"),
	(b"00000000010110000100001011010100", b"10010111111111001111000001011110"), -- -1.63458e-24 + 8.1055e-39 = -1.63458e-24
	(b"10100011101001100101000101100111", b"00000000000000000000000000000000"),
	(b"00000000011100110011010100111011", b"10100011101001100101000101100111"), -- -1.80322e-17 + 1.05802e-38 = -1.80322e-17
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001100101010001000111001", b"11111111100000000000000000000000"), -- -inf + -4.64997e-39 = -inf
	(b"10001100001010110101111000011100", b"00000000000000000000000000000000"),
	(b"10000000010010010111001100010101", b"10001100001010110101111000011101"), -- -1.32017e-31 + -6.74527e-39 = -1.32017e-31
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001111100101100101000110", b"01111111100000000000000000000000"), -- inf + -5.72583e-39 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100110100011111000000", b"10000000000100110100011111000000"), -- 0 + -1.77061e-39 = -1.77061e-39
	(b"01001000010001000000011110111101", b"00000000000000000000000000000000"),
	(b"10000000001111100110000001011011", b"01001000010001000000011110111101"), -- 200735 + -5.72837e-39 = 200735
	(b"10101000101111101110111101100001", b"00000000000000000000000000000000"),
	(b"00000000010000010110111011001111", b"10101000101111101110111101100001"), -- -2.11981e-14 + 6.00906e-39 = -2.11981e-14
	(b"11110010110000000101101011000000", b"00000000000000000000000000000000"),
	(b"10000000000010001000110011100011", b"11110010110000000101101011000000"), -- -7.61995e+30 + -7.85225e-40 = -7.61995e+30
	(b"10110010001000001100000000010010", b"00000000000000000000000000000000"),
	(b"00000000010010000000101110001011", b"10110010001000001100000000010010"), -- -9.3569e-09 + 6.6163e-39 = -9.3569e-09
	(b"01011100100011100101011101101001", b"00000000000000000000000000000000"),
	(b"10000000010010011101111001111010", b"01011100100011100101011101101001"), -- 3.20524e+17 + -6.7838e-39 = 3.20524e+17
	(b"00111001100001001001110001110100", b"00000000000000000000000000000000"),
	(b"10000000000100001001101110000010", b"00111001100001001001110001110100"), -- 0.000252936 + -1.52515e-39 = 0.000252936
	(b"00101011010111101000110001010110", b"00000000000000000000000000000000"),
	(b"00000000001111011011011000101001", b"00101011010111101000110001010110"), -- 7.9065e-13 + 5.66731e-39 = 7.9065e-13
	(b"00011001011100011110000100100011", b"00000000000000000000000000000000"),
	(b"00000000010110010000100010110010", b"00011001011100011110000100100011"), -- 1.25049e-23 + 8.17648e-39 = 1.25049e-23
	(b"10011001000011111001110101100000", b"00000000000000000000000000000000"),
	(b"10000000010110001101111000010001", b"10011001000011111001110101100000"), -- -7.42471e-24 + -8.16119e-39 = -7.42471e-24
	(b"01001111111101101010111010100111", b"00000000000000000000000000000000"),
	(b"10000000001101110101111000011111", b"01001111111101101010111010100111"), -- 8.27728e+09 + -5.08472e-39 = 8.27728e+09
	(b"11100101010010101111100001011101", b"00000000000000000000000000000000"),
	(b"10000000011100000111010110011100", b"11100101010010101111100001011101"), -- -5.99062e+22 + -1.03278e-38 = -5.99062e+22
	(b"00000000000000000000110100110000", b"00000000000000000000000000000000"),
	(b"10000000010001101100011100000000", b"10000000010001101011100111010000"), -- 4.73078e-42 + -6.49987e-39 = -6.49514e-39
	(b"10111000001100010011000100100100", b"00000000000000000000000000000000"),
	(b"10000000000000111101101001010011", b"10111000001100010011000100100100"), -- -4.22459e-05 + -3.53826e-40 = -4.22459e-05
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001100000110001101011011", b"11111111100000000000000000000000"), -- -inf + 4.44375e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011000010011110100010", b"11111111100000000000000000000000"), -- -inf + 9.93245e-39 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011111010100101011000110", b"11111111100000000000000000000000"), -- -inf + -1.15063e-38 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011100001100111110000110", b"01111111100000000000000000000000"), -- inf + -1.036e-38 = inf
	(b"10111000011100111101011111110000", b"00000000000000000000000000000000"),
	(b"00000000011001100111101100000011", b"10111000011100111101011111110000"), -- -5.81368e-05 + 9.41135e-39 = -5.81368e-05
	(b"11001011011011110000010111110001", b"00000000000000000000000000000000"),
	(b"00000000000000110111101110111011", b"11001011011011110000010111110001"), -- -1.56646e+07 + 3.19893e-40 = -1.56646e+07
	(b"00100100111000100011010100000101", b"00000000000000000000000000000000"),
	(b"00000000001001011100011111001010", b"00100100111000100011010100000101"), -- 9.81017e-17 + 3.46958e-39 = 9.81017e-17
	(b"00001010100000101111000111000000", b"00000000000000000000000000000000"),
	(b"10000000001010111110001111110010", b"00001010100000101111000110111101"), -- 1.26095e-32 + -4.0307e-39 = 1.26095e-32
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000011110010100010001001", b"11111111100000000000000000000000"), -- -inf + 1.39207e-39 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000010001011100110110110100", b"01111111100000000000000000000000"), -- inf + 6.41044e-39 = inf
	(b"11110101000100011111111011011011", b"00000000000000000000000000000000"),
	(b"00000000010101001011110011100011", b"11110101000100011111111011011011"), -- -1.85071e+32 + 7.78194e-39 = -1.85071e+32
	(b"11000111011100010011110110111010", b"00000000000000000000000000000000"),
	(b"10000000011000010011101010000011", b"11000111011100010011110110111010"), -- -61757.7 + -8.92903e-39 = -61757.7
	(b"01100010101001100001011101000100", b"00000000000000000000000000000000"),
	(b"10000000011111111001000011010001", b"01100010101001100001011101000100"), -- 1.53192e+21 + -1.17151e-38 = 1.53192e+21
	(b"10000000000000000000001000011000", b"00000000000000000000000000000000"),
	(b"00000000001100010001110000010010", b"00000000001100010001100111111010"), -- -7.51096e-43 + 4.51001e-39 = 4.50926e-39
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001110011100010110111011", b"01111111100000000000000000000000"), -- inf + 5.30556e-39 = inf
	(b"00000000000000000000101000001100", b"00000000000000000000000000000000"),
	(b"00000000001001110110000010011001", b"00000000001001110110101010100101"), -- 3.60414e-42 + 3.61624e-39 = 3.61984e-39
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011001100000111010010000", b"10000000011001100000111010010000"), -- 0 + -9.37244e-39 = -9.37244e-39
	(b"00101001100110110100111100010110", b"00000000000000000000000000000000"),
	(b"10000000001101110011011001000111", b"00101001100110110100111100010110"), -- 6.8971e-14 + -5.07042e-39 = 6.8971e-14
	(b"00110010100010011000101001010011", b"00000000000000000000000000000000"),
	(b"10000000000111110111100100010110", b"00110010100010011000101001010011"), -- 1.60118e-08 + -2.89034e-39 = 1.60118e-08
	(b"10111001010000111010011110101101", b"00000000000000000000000000000000"),
	(b"10000000011100100010010110011010", b"10111001010000111010011110101101"), -- -0.000186591 + -1.04827e-38 = -0.000186591
	(b"10000000000001011101110100010000", b"00000000000000000000000000000000"),
	(b"00000000000011111010101001100001", b"00000000000010011100110101010001"), -- -5.3848e-40 + 1.43865e-39 = 9.00173e-40
	(b"00000001100101100010100001010001", b"00000000000000000000000000000000"),
	(b"00000000011000000010010010101001", b"00000001101011100011000101111011"), -- 5.51591e-38 + 8.82936e-39 = 6.39885e-38
	(b"01010101100000010101100101001111", b"00000000000000000000000000000000"),
	(b"10000000001111000010111010000111", b"01010101100000010101100101001111"), -- 1.77776e+13 + -5.52682e-39 = 1.77776e+13
	(b"01010111111100110000001110110000", b"00000000000000000000000000000000"),
	(b"00000000011100110100110100110010", b"01010111111100110000001110110000"), -- 5.34394e+14 + 1.05888e-38 = 5.34394e+14
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000001101101010000011000011", b"11111111100000000000000000000000"), -- -inf + 5.01679e-39 = -inf
	(b"11010110000111100101110000001011", b"00000000000000000000000000000000"),
	(b"10000000001111010000110111010110", b"11010110000111100101110000001011"), -- -4.35295e+13 + -5.60693e-39 = -4.35295e+13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000101010010111000011011", b"01111111100000000000000000000000"), -- inf + 1.94508e-39 = inf
	(b"01110011000010100100100100100000", b"00000000000000000000000000000000"),
	(b"10000000011110001000110101100001", b"01110011000010100100100100100000"), -- 1.09561e+31 + -1.1071e-38 = 1.09561e+31
	(b"00100111100001001011110000000000", b"00000000000000000000000000000000"),
	(b"10000000011110000111101101010111", b"00100111100001001011110000000000"), -- 3.68412e-15 + -1.10645e-38 = 3.68412e-15
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001000010001010001110", b"00000000000001000010001010001110"), -- 0 + 3.79738e-40 = 3.79738e-40
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000011110010001000011010101", b"11111111100000000000000000000000"), -- -inf + -1.11181e-38 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000100010000100011111101", b"10000000000100010000100011111101"), -- 0 + -1.56443e-39 = -1.56443e-39
	(b"11011000100010111100010110001000", b"00000000000000000000000000000000"),
	(b"10000000000010000100001100110000", b"11011000100010111100010110001000"), -- -1.22944e+15 + -7.58786e-40 = -1.22944e+15
	(b"00101111011010100010000000010001", b"00000000000000000000000000000000"),
	(b"10000000001110111110110010011010", b"00101111011010100010000000010001"), -- 2.12936e-10 + -5.50317e-39 = 2.12936e-10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000011010100101110001100011", b"11111111100000000000000000000000"), -- -inf + 9.7677e-39 = -inf
	(b"11011001110101010001100000001100", b"00000000000000000000000000000000"),
	(b"10000000011111011101000100101011", b"11011001110101010001100000001100"), -- -7.49758e+15 + -1.15545e-38 = -7.49758e+15
	(b"10000001110110001001001000101110", b"00000000000000000000000000000000"),
	(b"00000000010001111011011100100011", b"10000001110001101010010001100101"), -- -7.95556e-38 + 6.58602e-39 = -7.29696e-38
	(b"11100000000010001010011100011110", b"00000000000000000000000000000000"),
	(b"10000000011111011110101000000111", b"11100000000010001010011100011110"), -- -3.93875e+19 + -1.15634e-38 = -3.93875e+19
	(b"00110000101111000000000101001010", b"00000000000000000000000000000000"),
	(b"00000000011111111011011100011001", b"00110000101111000000000101001010"), -- 1.36792e-09 + 1.17288e-38 = 1.36792e-09
	
	(b"00000000000110111110010000010011", b"00000000000000000000000000000000"),
	(b"10000000011000101111100010000000", b"10000000010001110001010001101101"), -- 2.56138e-39 + -9.08902e-39 = -6.52765e-39
	(b"00000000001010001011100001111000", b"00000000000000000000000000000000"),
	(b"00000000000010100111010001010011", b"00000000001100110010110011001011"), -- 3.73959e-39 + 9.60084e-40 = 4.69968e-39
	(b"10000000010100101011011110110100", b"00000000000000000000000000000000"),
	(b"00000000000010111111110010101100", b"10000000010001101011101100001000"), -- -7.59641e-39 + 1.10083e-39 = -6.49558e-39
	(b"00000000010110111011000001011010", b"00000000000000000000000000000000"),
	(b"10000000001001010010110000100101", b"00000000001101101000010000110101"), -- 8.42029e-39 + -3.41375e-39 = 5.00654e-39
	(b"00000000000110111011010000100001", b"00000000000000000000000000000000"),
	(b"00000000010001011011001011000001", b"00000000011000010110011011100010"), -- 2.54418e-39 + 6.40077e-39 = 8.94495e-39
	(b"10000000011011001010101111000100", b"00000000000000000000000000000000"),
	(b"00000000000011100010001000100111", b"10000000010111101000100110011101"), -- -9.97985e-39 + 1.29795e-39 = -8.6819e-39
	(b"10000000001110000001011000100000", b"00000000000000000000000000000000"),
	(b"10000000001100011000011011010011", b"10000000011010011001110011110011"), -- -5.15072e-39 + -4.54831e-39 = -9.69903e-39
	(b"10000000010011111000100111111011", b"00000000000000000000000000000000"),
	(b"00000000011111000010100100000011", b"00000000001011001001111100001000"), -- -7.3045e-39 + 1.14023e-38 = 4.09781e-39
	(b"00000000001101110001010000111101", b"00000000000000000000000000000000"),
	(b"10000000000001100101100000000011", b"00000000001100001011110000111010"), -- 5.05821e-39 + -5.82586e-40 = 4.47563e-39
	(b"10000000001101011110000111001110", b"00000000000000000000000000000000"),
	(b"00000000001000011110111101010110", b"10000000000100111111001001111000"), -- -4.94828e-39 + 3.11643e-39 = -1.83186e-39
	(b"10000000000011111100110101110111", b"00000000000000000000000000000000"),
	(b"00000000010011011100110010101110", b"00000000001111011111111100110111"), -- -1.45124e-39 + 7.14476e-39 = 5.69352e-39
	(b"10000000000011110110010000000011", b"00000000000000000000000000000000"),
	(b"10000000011000101011110110001001", b"10000000011100100010000110001100"), -- -1.41341e-39 + -9.06787e-39 = -1.04813e-38
	(b"10000000001100111111100001001100", b"00000000000000000000000000000000"),
	(b"10000000000101011101001110010110", b"10000000010010011100101111100010"), -- -4.77268e-39 + -2.00445e-39 = -6.77713e-39
	(b"10000000000111010001110011100001", b"00000000000000000000000000000000"),
	(b"10000000001011110110100010111001", b"10000000010011001000010110011010"), -- -2.67359e-39 + -4.35384e-39 = -7.02742e-39
	(b"10000000000101000010000110011101", b"00000000000000000000000000000000"),
	(b"00000000010110111001001000100100", b"00000000010001110111000010000111"), -- -1.84877e-39 + 8.40946e-39 = 6.56069e-39
	(b"00000000001110001011110100110110", b"00000000000000000000000000000000"),
	(b"00000000000110011000110110100101", b"00000000010100100100101011011011"), -- 5.21066e-39 + 2.3467e-39 = 7.55736e-39
	(b"00000000000010000100001010010000", b"00000000000000000000000000000000"),
	(b"00000000000100001001111100101110", b"00000000000110001110000110111110"), -- 7.58562e-40 + 1.52647e-39 = 2.28503e-39
	(b"10000000010001101001110001001010", b"00000000000000000000000000000000"),
	(b"00000000011100100011111100110011", b"00000000001010111010001011101001"), -- -6.48455e-39 + 1.04919e-38 = 4.00737e-39
	(b"00000000010000011001111000010000", b"00000000000000000000000000000000"),
	(b"10000000000011001010110011011110", b"00000000001101001111000100110010"), -- 6.02601e-39 + -1.16404e-39 = 4.86197e-39
	(b"10000000011110111011011001001100", b"00000000000000000000000000000000"),
	(b"10000000011010001101111001000101", b"10000000111001001001010010010001"), -- -1.13612e-38 + -9.63063e-39 = -2.09918e-38
	(b"10000000001000100111110001010110", b"00000000000000000000000000000000"),
	(b"00000000000100101010010110010110", b"10000000000011111101011011000000"), -- -3.16701e-39 + 1.71244e-39 = -1.45457e-39
	(b"10000000010011001110100110100100", b"00000000000000000000000000000000"),
	(b"00000000010000010110001110101010", b"10000000000010111000010111111010"), -- -7.06331e-39 + 6.00506e-39 = -1.05825e-39
	(b"00000000000001100100011000100111", b"00000000000000000000000000000000"),
	(b"00000000001000001110101100010100", b"00000000001001110011000100111011"), -- 5.76179e-40 + 3.02307e-39 = 3.59924e-39
	(b"00000000000110101000010100110100", b"00000000000000000000000000000000"),
	(b"10000000001010010011001001101101", b"10000000000011101010110100111001"), -- 2.43551e-39 + -3.78334e-39 = -1.34784e-39
	(b"10000000010001000100010001111101", b"00000000000000000000000000000000"),
	(b"00000000011101101010101111011010", b"00000000001100100110011101011101"), -- -6.26938e-39 + 1.08982e-38 = 4.62885e-39
	(b"00000000001010111001111101111010", b"00000000000000000000000000000000"),
	(b"10000000011010000000011010011010", b"10000000001111000110011100100000"), -- 4.00614e-39 + -9.55326e-39 = -5.54712e-39
	(b"00000000010110100011110110000101", b"00000000000000000000000000000000"),
	(b"10000000011001010101001000001111", b"10000000000010110001010010001010"), -- 8.28726e-39 + -9.30482e-39 = -1.01756e-39
	(b"10000000001110110011001100101000", b"00000000000000000000000000000000"),
	(b"00000000011111111001100111000111", b"00000000010001000110011010011111"), -- -5.43665e-39 + 1.17183e-38 = 6.28163e-39
	(b"10000000010100110100110101011110", b"00000000000000000000000000000000"),
	(b"10000000000100000110010110010100", b"10000000011000111011001011110010"), -- -7.6501e-39 + -1.50581e-39 = -9.15591e-39
	(b"00000000001100000001000010111010", b"00000000000000000000000000000000"),
	(b"00000000001100011101010101111010", b"00000000011000011110011000110100"), -- 4.4141e-39 + 4.57652e-39 = 8.99062e-39
	(b"00000000010101001110111111010101", b"00000000000000000000000000000000"),
	(b"00000000001110001011011010101111", b"00000000100011011010011010000100"), -- 7.80022e-39 + 5.20832e-39 = 1.30085e-38
	(b"00000000011101110101110001111101", b"00000000000000000000000000000000"),
	(b"00000000001100000100001101101111", b"00000000101001111001111111101100"), -- 1.09616e-38 + 4.43229e-39 = 1.53939e-38
	(b"10000000010010101001101001011110", b"00000000000000000000000000000000"),
	(b"10000000011111001101110100011010", b"10000000110001110111011101111000"), -- -6.8512e-39 + -1.14669e-38 = -1.83181e-38
	(b"00000000000110000011100011101001", b"00000000000000000000000000000000"),
	(b"10000000001100010100101101110111", b"10000000000110010001001010001110"), -- 2.22447e-39 + -4.52701e-39 = -2.30254e-39
	(b"00000000000110110000101111110101", b"00000000000000000000000000000000"),
	(b"10000000010000101110011101110100", b"10000000001001111101101101111111"), -- 2.48385e-39 + -6.14417e-39 = -3.66032e-39
	(b"10000000001110000110001111001110", b"00000000000000000000000000000000"),
	(b"10000000001100110101111000100111", b"10000000011010111100000111110101"), -- -5.17859e-39 + -4.71739e-39 = -9.89598e-39
	(b"00000000011010110110010100100100", b"00000000000000000000000000000000"),
	(b"00000000000111101111001010100111", b"00000000100010100101011111001011"), -- 9.86268e-39 + 2.84211e-39 = 1.27048e-38
	(b"00000000000011001100011111011001", b"00000000000000000000000000000000"),
	(b"10000000001110001111101110111011", b"10000000001011000011001111100010"), -- 1.17372e-39 + -5.23309e-39 = -4.05937e-39
	(b"00000000001100111111101010110110", b"00000000000000000000000000000000"),
	(b"00000000011011000001101011001101", b"00000000101000000001010110000011"), -- 4.77355e-39 + 9.92785e-39 = 1.47014e-38
	(b"10000000010001101111001101011101", b"00000000000000000000000000000000"),
	(b"00000000010010110011101100011010", b"00000000000001000100011110111101"), -- -6.51579e-39 + 6.90886e-39 = 3.93077e-40
	(b"10000000010111111101001110101110", b"00000000000000000000000000000000"),
	(b"00000000010111101011000000100111", b"10000000000000010010001110000111"), -- -8.80031e-39 + 8.69573e-39 = -1.0458e-40
	(b"00000000001001010010001011011100", b"00000000000000000000000000000000"),
	(b"00000000000111010000100111100110", b"00000000010000100010110011000010"), -- 3.41042e-39 + 2.66678e-39 = 6.0772e-39
	(b"00000000001000011001011100110010", b"00000000000000000000000000000000"),
	(b"10000000011111010000010100000100", b"10000000010110110110110111010010"), -- 3.08481e-39 + -1.14812e-38 = -8.39643e-39
	(b"10000000011101100011100011010101", b"00000000000000000000000000000000"),
	(b"10000000011111101101001110111011", b"10000000111101010000110010010000"), -- -1.0857e-38 + -1.16472e-38 = -2.25042e-38
	(b"00000000000000011001100110011000", b"00000000000000000000000000000000"),
	(b"00000000010100101100110101111011", b"00000000010101000110011100010011"), -- 1.46935e-40 + 7.60422e-39 = 7.75116e-39
	(b"00000000000110011111011010110011", b"00000000000000000000000000000000"),
	(b"10000000010100000000011110101111", b"10000000001101100001000011111100"), -- 2.38439e-39 + -7.3496e-39 = -4.96521e-39
	(b"00000000010110000010011100001110", b"00000000000000000000000000000000"),
	(b"00000000001011011000000111111000", b"00000000100001011010100100000110"), -- 8.09553e-39 + 4.17922e-39 = 1.22748e-38
	(b"00000000001100000011110001111011", b"00000000000000000000000000000000"),
	(b"10000000011000001101110111110100", b"10000000001100001010000101111001"), -- 4.4298e-39 + -8.89583e-39 = -4.46603e-39
	(b"10000000010101000111000000110111", b"00000000000000000000000000000000"),
	(b"00000000011100101001010110011101", b"00000000000111100010010101100110"), -- -7.75444e-39 + 1.05229e-38 = 2.76848e-39
	(b"00000000001100001000000100100110", b"00000000000000000000000000000000"),
	(b"00000000001100011000010100111110", b"00000000011000100000011001100100"), -- 4.45443e-39 + 4.54774e-39 = 9.00217e-39
	(b"00000000001001011101010110100101", b"00000000000000000000000000000000"),
	(b"10000000000110111110101011101001", b"00000000000010011110101010111100"), -- 3.47455e-39 + -2.56383e-39 = 9.10726e-40
	(b"00000000010011011101101101010001", b"00000000000000000000000000000000"),
	(b"10000000011110101001010000101011", b"10000000001011001011100011011010"), -- 7.15001e-39 + -1.12571e-38 = -4.10707e-39
	(b"00000000011000001000100001100111", b"00000000000000000000000000000000"),
	(b"00000000010100000001110101000100", b"00000000101100001010010110101011"), -- 8.86514e-39 + 7.35734e-39 = 1.62225e-38
	(b"00000000000011011110111110101100", b"00000000000000000000000000000000"),
	(b"00000000001111010101110010000010", b"00000000010010110100110000101110"), -- 1.27984e-39 + 5.63515e-39 = 6.91499e-39
	(b"10000000010011100101011010010001", b"00000000000000000000000000000000"),
	(b"00000000010001011010011100110011", b"10000000000010001010111101011110"), -- -7.19422e-39 + 6.39663e-39 = -7.97594e-40
	(b"00000000011111011100101000110101", b"00000000000000000000000000000000"),
	(b"00000000001101111101100101101000", b"00000000101101011010001110011101"), -- 1.1552e-38 + 5.12894e-39 = 1.66809e-38
	(b"00000000000010111100001010010000", b"00000000000000000000000000000000"),
	(b"00000000001000000001000010010000", b"00000000001010111101001100100000"), -- 1.07999e-39 + 2.94468e-39 = 4.02466e-39
	(b"00000000000111110100100010000111", b"00000000000000000000000000000000"),
	(b"10000000011110010110001000010110", b"10000000010110100001100110001111"), -- 2.87292e-39 + -1.11473e-38 = -8.27436e-39
	(b"10000000010001010110101100010100", b"00000000000000000000000000000000"),
	(b"00000000011011100010110100101100", b"00000000001010001100001000011000"), -- -6.37506e-39 + 1.01181e-38 = 3.74305e-39
	(b"00000000001001110111101011111000", b"00000000000000000000000000000000"),
	(b"00000000011100010100010110111010", b"00000000100110001100000010110010"), -- 3.6257e-39 + 1.04024e-38 = 1.40281e-38
	(b"10000000010110011000110111100011", b"00000000000000000000000000000000"),
	(b"00000000001110100010011010011001", b"10000000000111110110011101001010"), -- -8.22426e-39 + 5.34031e-39 = -2.88395e-39
	(b"00000000001000011101010010010110", b"00000000000000000000000000000000"),
	(b"10000000001001010101001011111011", b"10000000000000110111111001100101"), -- 3.10683e-39 + -3.42768e-39 = -3.20848e-40
	(b"10000000011010000101111110000010", b"00000000000000000000000000000000"),
	(b"10000000001001000100011111100100", b"10000000100011001010011101100110"), -- -9.58515e-39 + -3.33187e-39 = -1.2917e-38
	(b"10000000011000100001101010110001", b"00000000000000000000000000000000"),
	(b"00000000011001101010000011010011", b"00000000000001001000011000100010"), -- -9.00945e-39 + 9.42491e-39 = 4.1546e-40
	(b"10000000000101111100100000000001", b"00000000000000000000000000000000"),
	(b"10000000011000110001100010101011", b"10000000011110101110000010101100"), -- -2.18396e-39 + -9.10056e-39 = -1.12845e-38
	(b"00000000001110111101100001100000", b"00000000000000000000000000000000"),
	(b"10000000001011111101011001010011", b"00000000000011000000001000001101"), -- 5.49591e-39 + -4.39315e-39 = 1.10276e-39
	(b"00000000000001011111010101110100", b"00000000000000000000000000000000"),
	(b"00000000011111011101100110100100", b"00000000100000111100111100011000"), -- 5.47229e-40 + 1.15575e-38 = 1.21047e-38
	(b"00000000010000011111010101010010", b"00000000000000000000000000000000"),
	(b"10000000000011001010011011000111", b"00000000001101010100111010001011"), -- 6.05731e-39 + -1.16185e-39 = 4.89546e-39
	(b"00000000010001100100111111111101", b"00000000000000000000000000000000"),
	(b"00000000011111010110100000011101", b"00000000110000111011100000011010"), -- 6.45718e-39 + 1.15168e-38 = 1.7974e-38
	(b"00000000001001111010011011001111", b"00000000000000000000000000000000"),
	(b"10000000000010110110011111000000", b"00000000000111000011111100001111"), -- 3.64142e-39 + -1.04741e-39 = 2.59402e-39
	(b"10000000011011001100001001100100", b"00000000000000000000000000000000"),
	(b"10000000000001111000111000001000", b"10000000011101000101000001101100"), -- -9.98797e-39 + -6.938e-40 = -1.06818e-38
	(b"00000000010000000000010101111101", b"00000000000000000000000000000000"),
	(b"10000000011101111100101111111100", b"10000000001101111100011001111111"), -- 5.87944e-39 + -1.10016e-38 = -5.12216e-39
	(b"00000000000000011100010001111011", b"00000000000000000000000000000000"),
	(b"10000000011010101101011001010010", b"10000000011010010001000111010111"), -- 1.62319e-40 + -9.81145e-39 = -9.64913e-39
	(b"10000000011000000111010110001010", b"00000000000000000000000000000000"),
	(b"10000000000110001101000101010100", b"10000000011110010100011011011110"), -- -8.85837e-39 + -2.27914e-39 = -1.11375e-38
	(b"10000000011011110111100101111101", b"00000000000000000000000000000000"),
	(b"00000000001000000100110011010100", b"10000000010011110010110010101001"), -- -1.02373e-38 + 2.9663e-39 = -7.27103e-39
	(b"10000000001010101010001010000110", b"00000000000000000000000000000000"),
	(b"00000000010100111011000000101100", b"00000000001010010000110110100110"), -- -3.91539e-39 + 7.68554e-39 = 3.77015e-39
	(b"00000000010100100010001001111110", b"00000000000000000000000000000000"),
	(b"00000000011011011001101101001100", b"00000000101111111011110111001010"), -- 7.54288e-39 + 1.00658e-38 = 1.76087e-38
	(b"00000000011111010111101000101110", b"00000000000000000000000000000000"),
	(b"10000000001100110100000111111001", b"00000000010010100011100000110101"), -- 1.15233e-38 + -4.70728e-39 = 6.81599e-39
	(b"00000000010000110011111000001000", b"00000000000000000000000000000000"),
	(b"00000000011110101011010000001111", b"00000000101111011111001000010111"), -- 6.17523e-39 + 1.12685e-38 = 1.74438e-38
	(b"00000000010000111000011010011110", b"00000000000000000000000000000000"),
	(b"10000000011010010001111011110110", b"10000000001001011001100001011000"), -- 6.20127e-39 + -9.65383e-39 = -3.45256e-39
	(b"00000000000001011100010000011101", b"00000000000000000000000000000000"),
	(b"00000000010101010010111110110111", b"00000000010110101111001111010100"), -- 5.2953e-40 + 7.82313e-39 = 8.35266e-39
	(b"00000000000011111011110001000101", b"00000000000000000000000000000000"),
	(b"00000000011110010100110011010011", b"00000000100010010000100100011000"), -- 1.44507e-39 + 1.11397e-38 = 1.25847e-38
	(b"00000000000100000010101011101101", b"00000000000000000000000000000000"),
	(b"10000000011110100101010011011110", b"10000000011010100010100111110001"), -- 1.48477e-39 + -1.12344e-38 = -9.74961e-39
	(b"00000000000101011100101011110000", b"00000000000000000000000000000000"),
	(b"10000000011101001101101000001111", b"10000000010111110000111100011111"), -- 2.00135e-39 + -1.07311e-38 = -8.7298e-39
	(b"00000000010000001101100000010100", b"00000000000000000000000000000000"),
	(b"10000000011101010110101011000111", b"10000000001101001001001010110011"), -- 5.95499e-39 + -1.07831e-38 = -4.82807e-39
	(b"00000000010011111100011000100011", b"00000000000000000000000000000000"),
	(b"00000000000110110001110011010100", b"00000000011010101110001011110111"), -- 7.32608e-39 + 2.4899e-39 = 9.81598e-39
	(b"00000000000101110111000101000001", b"00000000000000000000000000000000"),
	(b"00000000010110001100001100100101", b"00000000011100000011010001100110"), -- 2.15284e-39 + 8.15153e-39 = 1.03044e-38
	(b"10000000000011010001100100110000", b"00000000000000000000000000000000"),
	(b"10000000011110011111001101101000", b"10000000100001110000110010011000"), -- -1.2029e-39 + -1.11994e-38 = -1.24023e-38
	(b"00000000000000101101111111101001", b"00000000000000000000000000000000"),
	(b"10000000001101111100110000101101", b"10000000001101001110110001000100"), -- 2.63995e-40 + -5.1242e-39 = -4.8602e-39
	(b"10000000010000100010001100101010", b"00000000000000000000000000000000"),
	(b"10000000001101101001000111101110", b"10000000011110001011010100011000"), -- -6.07376e-39 + -5.01147e-39 = -1.10852e-38
	(b"00000000010011111011100000100011", b"00000000000000000000000000000000"),
	(b"10000000011011101000100101110010", b"10000000000111101101000101001111"), -- 7.32106e-39 + -1.01512e-38 = -2.83015e-39
	(b"00000000001011011000111000101000", b"00000000000000000000000000000000"),
	(b"00000000010110111110000100011100", b"00000000100010010110111101000100"), -- 4.18359e-39 + 8.43778e-39 = 1.26214e-38
	(b"10000000011111100100011011011001", b"00000000000000000000000000000000"),
	(b"10000000011001011111000111111111", b"10000000111001000011100011011000"), -- -1.15967e-38 + -9.3622e-39 = -2.09589e-38
	(b"10000000011101111010010111000101", b"00000000000000000000000000000000"),
	(b"00000000000000011011101101000011", b"10000000011101011110101010000010"), -- -1.09879e-38 + 1.59012e-40 = -1.08289e-38
	(b"00000000001101010111001011001110", b"00000000000000000000000000000000"),
	(b"10000000000000101000001110101111", b"00000000001100101110111100011111"), -- 4.90847e-39 + -2.3091e-40 = 4.67756e-39
	(b"10000000001111101111101001010010", b"00000000000000000000000000000000"),
	(b"10000000010101101100000111000011", b"10000000100101011011110000010101"), -- -5.7836e-39 + -7.96736e-39 = -1.3751e-38
	(b"10000000000001000111000110101000", b"00000000000000000000000000000000"),
	(b"00000000000110001101010100101011", b"00000000000101000110001110000011"), -- -4.08114e-40 + 2.28052e-39 = 1.87241e-39
	(b"00000000011010011011100001000100", b"00000000000000000000000000000000"),
	(b"00000000000001101011101000101100", b"00000000011100000111001001110000"), -- 9.70883e-39 + 6.17799e-40 = 1.03266e-38
	(b"00000000010010100111010101000110", b"00000000000000000000000000000000"),
	(b"10000000000110001001100101011011", b"00000000001100011101101111101011"), -- 6.8379e-39 + -2.25907e-39 = 4.57883e-39
	(b"00000000001011110110100000010101", b"00000000000000000000000000000000"),
	(b"10000000001001011000110101000001", b"00000000000010011101101011010100"), -- 4.35361e-39 + -3.44859e-39 = 9.0502e-40
	(b"00000000000011000101001101100100", b"00000000000000000000000000000000"),
	(b"10000000010111111010011010010001", b"10000000010100110101001100101101"), -- 1.13194e-39 + -8.78412e-39 = -7.65218e-39
	(b"10000000011010000110101001111101", b"00000000000000000000000000000000"),
	(b"10000000010111111011011101011100", b"10000000110010000010000111011001"), -- -9.58909e-39 + -8.79015e-39 = -1.83792e-38
	(b"10000000011011000011111010001111", b"00000000000000000000000000000000"),
	(b"10000000011101111101101011010111", b"10000000111001000001100101100110"), -- -9.94068e-39 + -1.10069e-38 = -2.09476e-38
	(b"10000000000110110010011010110100", b"00000000000000000000000000000000"),
	(b"00000000000011111101111001111011", b"10000000000010110100100000111001"), -- -2.49344e-39 + 1.45734e-39 = -1.0361e-39
	(b"10000000011100010010101100111011", b"00000000000000000000000000000000"),
	(b"00000000001001001000110001001101", b"10000000010011001001111011101110"), -- -1.03929e-38 + 3.35641e-39 = -7.03651e-39
	(b"10000000010111100001000000001011", b"00000000000000000000000000000000"),
	(b"10000000010101010010100011001000", b"10000000101100110011100011010011"), -- -8.63829e-39 + -7.82065e-39 = -1.64589e-38
	(b"00000000010101000101110101000011", b"00000000000000000000000000000000"),
	(b"00000000010111100100101110000010", b"00000000101100101010100011000101"), -- 7.74764e-39 + 8.65962e-39 = 1.64073e-38
	(b"00000000011001001110101010011111", b"00000000000000000000000000000000"),
	(b"10000000010000000111100101100001", b"00000000001001000111000100111110"), -- 9.26772e-39 + -5.92101e-39 = 3.3467e-39
	(b"10000000001101000100101000110101", b"00000000000000000000000000000000"),
	(b"10000000011100001110101100001001", b"10000000101001010011010100111110"), -- -4.80207e-39 + -1.03699e-38 = -1.5172e-38
	(b"00000000001110000100101101100101", b"00000000000000000000000000000000"),
	(b"00000000011110101001110001011110", b"00000000101100101110011111000011"), -- 5.16983e-39 + 1.126e-38 = 1.64299e-38
	(b"00000000001010100000001101010011", b"00000000000000000000000000000000"),
	(b"10000000011011110110011000110100", b"10000000010001010110001011100001"), -- 3.85828e-39 + -1.02304e-38 = -6.37212e-39
	(b"00000000010010001100110110000001", b"00000000000000000000000000000000"),
	(b"00000000000110001101001111100000", b"00000000011000011010000101100001"), -- 6.68588e-39 + 2.28006e-39 = 8.96593e-39
	(b"00000000011011110000000100100111", b"00000000000000000000000000000000"),
	(b"00000000010000010001001010101101", b"00000000101100000001001111010100"), -- 1.01942e-38 + 5.97601e-39 = 1.61702e-38
	(b"10000000010011011000010010001111", b"00000000000000000000000000000000"),
	(b"00000000001011001111000000000001", b"10000000001000001001010010001110"), -- -7.11889e-39 + 4.12686e-39 = -2.99203e-39
	(b"10000000001011001011011011000000", b"00000000000000000000000000000000"),
	(b"10000000010100101010011001100011", b"10000000011111110101110100100011"), -- -4.10632e-39 + -7.5902e-39 = -1.16965e-38
	(b"00000000001000010001001101111110", b"00000000000000000000000000000000"),
	(b"00000000011010100100111000000011", b"00000000100010110110000110000001"), -- 3.03756e-39 + 9.76255e-39 = 1.28001e-38
	(b"10000000000110110110011111101100", b"00000000000000000000000000000000"),
	(b"10000000011011110110000000000010", b"10000000100010101100011111101110"), -- -2.51684e-39 + -1.02282e-38 = -1.2745e-38
	(b"10000000000011111110100100000110", b"00000000000000000000000000000000"),
	(b"00000000010010111010101101010100", b"00000000001110111100001001001110"), -- -1.46113e-39 + 6.94912e-39 = 5.488e-39
	(b"10000000011101000110011111011100", b"00000000000000000000000000000000"),
	(b"10000000011011001100100000100111", b"10000000111000010011000000000011"), -- -1.06902e-38 + -9.99003e-39 = -2.06802e-38
	(b"00000000010111100001011000110101", b"00000000000000000000000000000000"),
	(b"00000000011111001110101110011011", b"00000000110110110000000111010000"), -- 8.6405e-39 + 1.14721e-38 = 2.01126e-38
	(b"00000000000000010101100001110111", b"00000000000000000000000000000000"),
	(b"00000000010100010110011110100101", b"00000000010100101100000000011100"), -- 1.23571e-40 + 7.47586e-39 = 7.59943e-39
	(b"10000000000100101000001000111010", b"00000000000000000000000000000000"),
	(b"10000000010010011110101010111110", b"10000000010111000110110011111000"), -- -1.69976e-39 + -6.7882e-39 = -8.48796e-39
	(b"00000000001011001000101110000100", b"00000000000000000000000000000000"),
	(b"10000000001101010100111101110111", b"10000000000010001100001111110011"), -- 4.09081e-39 + -4.89579e-39 = -8.04977e-40
	(b"00000000000010101101011010010111", b"00000000000000000000000000000000"),
	(b"10000000000000000011011001110001", b"00000000000010101010000000100110"), -- 9.95335e-40 + -1.95299e-41 = 9.75805e-40
	(b"00000000011101100000001010110110", b"00000000000000000000000000000000"),
	(b"00000000010100011100101001011011", b"00000000110001111100110100010001"), -- 1.08376e-38 + 7.51127e-39 = 1.83488e-38
	(b"00000000001010101101110110100000", b"00000000000000000000000000000000"),
	(b"00000000000101110010010001110101", b"00000000010000100000001000010101"), -- 3.93659e-39 + 2.12529e-39 = 6.06189e-39
	(b"00000000000000101010010011101010", b"00000000000000000000000000000000"),
	(b"10000000011101100110111111111101", b"10000000011100111100101100010011"), -- 2.42831e-40 + -1.08768e-38 = -1.06339e-38
	(b"10000000010101010010011100111111", b"00000000000000000000000000000000"),
	(b"10000000010100010010010111001100", b"10000000101001100100110100001011"), -- -7.8201e-39 + -7.45223e-39 = -1.52723e-38
	(b"10000000000000101000100100101101", b"00000000000000000000000000000000"),
	(b"00000000010100011101110000001101", b"00000000010011110101001011100000"), -- -2.3288e-40 + 7.51761e-39 = 7.28473e-39
	(b"00000000000110000101011000010100", b"00000000000000000000000000000000"),
	(b"00000000010000101011111110111000", b"00000000010110110001010111001100"), -- 2.23493e-39 + 6.12992e-39 = 8.36485e-39
	(b"00000000010111000000111101100010", b"00000000000000000000000000000000"),
	(b"00000000010100101011111101010011", b"00000000101011101100111010110101"), -- 8.45438e-39 + 7.59914e-39 = 1.60535e-38
	(b"10000000010110100101100100001111", b"00000000000000000000000000000000"),
	(b"10000000011010011011110110011001", b"10000000110001000001011010101000"), -- -8.29714e-39 + -9.71074e-39 = -1.80079e-38
	(b"00000000011101001111110110000100", b"00000000000000000000000000000000"),
	(b"00000000001001110101100111100010", b"00000000100111000101011101100110"), -- 1.07439e-38 + 3.61383e-39 = 1.43577e-38
	(b"10000000011111100110000111100110", b"00000000000000000000000000000000"),
	(b"10000000001011001101101110101001", b"10000000101010110011110110001111"), -- -1.16064e-38 + -4.11956e-39 = -1.5726e-38
	(b"10000000010001001101110110001001", b"00000000000000000000000000000000"),
	(b"00000000001101111011010010001000", b"10000000000011010010100100000001"), -- -6.32429e-39 + 5.11571e-39 = -1.20857e-39
	(b"00000000001000011110110110010010", b"00000000000000000000000000000000"),
	(b"00000000000101011001010110001101", b"00000000001101111000001100011111"), -- 3.1158e-39 + 1.98219e-39 = 5.09799e-39
	(b"10000000010111111001011010010110", b"00000000000000000000000000000000"),
	(b"10000000011010110011011000011101", b"10000000110010101100110010110011"), -- -8.77839e-39 + -9.84581e-39 = -1.86242e-38
	(b"00000000000001010001110001100000", b"00000000000000000000000000000000"),
	(b"00000000001010111001001001111001", b"00000000001100001010111011011001"), -- 4.69357e-40 + 4.00147e-39 = 4.47083e-39
	(b"10000000010011011100000101100000", b"00000000000000000000000000000000"),
	(b"10000000000111010111100100010011", b"10000000011010110011101001110011"), -- -7.1407e-39 + -2.70666e-39 = -9.84737e-39
	(b"00000000011000010001111110000001", b"00000000000000000000000000000000"),
	(b"10000000010101010111011101111100", b"00000000000010111010100000000101"), -- 8.91934e-39 + -7.84888e-39 = 1.07046e-39
	(b"10000000010100100000000000101111", b"00000000000000000000000000000000"),
	(b"10000000001010111101011000110010", b"10000000011111011101011001100001"), -- -7.53058e-39 + -4.02577e-39 = -1.15563e-38
	(b"00000000010111111010110000011010", b"00000000000000000000000000000000"),
	(b"00000000001001000001110010100110", b"00000000100000111100100011000000"), -- 8.78611e-39 + 3.31635e-39 = 1.21025e-38
	(b"10000000001110111011101011110011", b"00000000000000000000000000000000"),
	(b"00000000001001000101110001001010", b"10000000000101110101111010101001"), -- -5.48536e-39 + 3.33918e-39 = -2.14617e-39
	(b"00000000000011011111110000011010", b"00000000000000000000000000000000"),
	(b"00000000001000100010011010111111", b"00000000001100000010001011011001"), -- 1.2843e-39 + 3.13631e-39 = 4.4206e-39
	(b"00000000000101111110110111011011", b"00000000000000000000000000000000"),
	(b"00000000001110000000110011000001", b"00000000010011111111101010011100"), -- 2.19754e-39 + 5.14736e-39 = 7.34491e-39
	(b"00000000000100000101000011010111", b"00000000000000000000000000000000"),
	(b"10000000011011101100011101101011", b"10000000010111100111011010010100"), -- 1.49837e-39 + -1.01734e-38 = -8.67507e-39
	(b"00000000001111101001101110011100", b"00000000000000000000000000000000"),
	(b"00000000000010101000111010100110", b"00000000010010010010101001000010"), -- 5.74962e-39 + 9.69528e-40 = 6.71915e-39
	(b"00000000010010001010101011100011", b"00000000000000000000000000000000"),
	(b"10000000001001100111010011010111", b"00000000001000100011011000001100"), -- 6.67346e-39 + -3.53166e-39 = 3.1418e-39
	(b"10000000001111000001111011000010", b"00000000000000000000000000000000"),
	(b"00000000010110000011010010100100", b"00000000000111000001010111100010"), -- -5.52116e-39 + 8.10041e-39 = 2.57924e-39
	(b"00000000000011001101111100000000", b"00000000000000000000000000000000"),
	(b"10000000011000100110011111111001", b"10000000010101011000100011111001"), -- 1.18202e-39 + -9.03718e-39 = -7.85515e-39
	(b"10000000001010110011000101010001", b"00000000000000000000000000000000"),
	(b"00000000011111101111111000001100", b"00000000010100111100110010111011"), -- -3.96662e-39 + 1.16624e-38 = 7.69579e-39
	(b"10000000000110001100010100001101", b"00000000000000000000000000000000"),
	(b"10000000011010010000000010010000", b"10000000100000011100010110011101"), -- -2.27474e-39 + -9.64293e-39 = -1.19177e-38
	(b"10000000001101010001111111010110", b"00000000000000000000000000000000"),
	(b"10000000000001101100010110000110", b"10000000001110111110010101011100"), -- -4.8787e-39 + -6.21871e-40 = -5.50057e-39
	(b"00000000001010100111100000110011", b"00000000000000000000000000000000"),
	(b"00000000011011100100110000011111", b"00000000100110001100010001010010"), -- 3.90021e-39 + 1.01292e-38 = 1.40294e-38
	(b"00000000011100100010110110111100", b"00000000000000000000000000000000"),
	(b"10000000001010101110000001011110", b"00000000010001110100110101011110"), -- 1.04857e-38 + -3.93758e-39 = 6.54807e-39
	(b"10000000011010110010010101110011", b"00000000000000000000000000000000"),
	(b"10000000000100000011001001111001", b"10000000011110110101011111101100"), -- -9.83983e-39 + -1.48747e-39 = -1.13273e-38
	(b"00000000001100011011111001000101", b"00000000000000000000000000000000"),
	(b"10000000010001101100111011011100", b"10000000000101010001000010010111"), -- 4.5682e-39 + -6.50269e-39 = -1.9345e-39
	(b"10000000001000100001101101110011", b"00000000000000000000000000000000"),
	(b"10000000010100111100100111001000", b"10000000011101011110010100111011"), -- -3.13225e-39 + -7.69473e-39 = -1.0827e-38
	(b"00000000000111010100111100000111", b"00000000000000000000000000000000"),
	(b"00000000011000010111010000111011", b"00000000011111101100001101000010"), -- 2.69158e-39 + 8.94974e-39 = 1.16413e-38
	(b"00000000001011110101111111111001", b"00000000000000000000000000000000"),
	(b"10000000010001101110100010110011", b"10000000000101111000100010111010"), -- 4.3507e-39 + -6.51196e-39 = -2.16126e-39
	(b"00000000000110101111010111111110", b"00000000000000000000000000000000"),
	(b"10000000010011001010000111100111", b"10000000001100011010101111101001"), -- 2.47597e-39 + -7.03758e-39 = -4.56161e-39
	(b"00000000011100001001000101010110", b"00000000000000000000000000000000"),
	(b"10000000010000001111001111011011", b"00000000001011111001110101111011"), -- 1.03377e-38 + -5.96495e-39 = 4.37276e-39
	(b"00000000011101001001101101000001", b"00000000000000000000000000000000"),
	(b"10000000001110111101001100101001", b"00000000001110001100100000011000"), -- 1.07086e-38 + -5.49404e-39 = 5.21457e-39
	(b"00000000000001001001110001000101", b"00000000000000000000000000000000"),
	(b"10000000010111101101000010111110", b"10000000010110100011010001111001"), -- 4.23401e-40 + -8.70742e-39 = -8.28402e-39
	(b"10000000010111011010110101011111", b"00000000000000000000000000000000"),
	(b"10000000001010010010111010100011", b"10000000100001101101110000000010"), -- -8.60289e-39 + -3.78199e-39 = -1.23849e-38
	(b"10000000001001111111000100101010", b"00000000000000000000000000000000"),
	(b"10000000010101001111101010100100", b"10000000011111001110101111001110"), -- -3.6681e-39 + -7.80409e-39 = -1.14722e-38
	(b"00000000000100000000101010000111", b"00000000000000000000000000000000"),
	(b"00000000001010101011000001101111", b"00000000001110101011101011110110"), -- 1.47314e-39 + 3.92038e-39 = 5.39353e-39
	(b"00000000010101010010001001110111", b"00000000000000000000000000000000"),
	(b"00000000001001000000101011110101", b"00000000011110010010110101101100"), -- 7.81838e-39 + 3.31001e-39 = 1.11284e-38
	(b"00000000001000000001111001110110", b"00000000000000000000000000000000"),
	(b"10000000010111010101011010101000", b"10000000001111010011100000110010"), -- 2.94966e-39 + -8.57179e-39 = -5.62212e-39
	(b"00000000000100100101100101111111", b"00000000000000000000000000000000"),
	(b"00000000011000110010101001011011", b"00000000011101011000001111011010"), -- 1.68514e-39 + 9.10691e-39 = 1.07921e-38
	(b"10000000001110101110111011001110", b"00000000000000000000000000000000"),
	(b"10000000000100010101000010110110", b"10000000010011000011111110000100"), -- -5.41213e-39 + -1.59016e-39 = -7.00228e-39
	(b"00000000000010011111010110000101", b"00000000000000000000000000000000"),
	(b"10000000011011000110011100001000", b"10000000011000100111000110000011"), -- 9.14595e-40 + -9.95519e-39 = -9.0406e-39
	(b"10000000001000011101111010111010", b"00000000000000000000000000000000"),
	(b"00000000000101011100100110011010", b"10000000000011000001010100100000"), -- -3.11047e-39 + 2.00087e-39 = -1.1096e-39
	(b"10000000010000110110010010101100", b"00000000000000000000000000000000"),
	(b"10000000010111101011011010101011", b"10000000101000100001101101010111"), -- -6.18909e-39 + -8.69807e-39 = -1.48872e-38
	(b"00000000000010010110001100111011", b"00000000000000000000000000000000"),
	(b"00000000011111111011000101100000", b"00000000100010010001010010011011"), -- 8.62117e-40 + 1.17267e-38 = 1.25889e-38
	(b"00000000010100010111111010110000", b"00000000000000000000000000000000"),
	(b"10000000001101110001101000001001", b"00000000000110100110010010100111"), -- 7.48412e-39 + -5.06029e-39 = 2.42383e-39
	(b"10000000010101101110101110000101", b"00000000000000000000000000000000"),
	(b"10000000011101001011110011011110", b"10000000110010111010100001100011"), -- -7.98234e-39 + -1.07207e-38 = -1.8703e-38
	(b"00000000011111010001100101110110", b"00000000000000000000000000000000"),
	(b"00000000000000111100110000001001", b"00000000100000001110010101111111"), -- 1.14886e-38 + 3.48701e-40 = 1.18373e-38
	(b"10000000000010011011000000100110", b"00000000000000000000000000000000"),
	(b"10000000001011101001001110001110", b"10000000001110000100001110110100"), -- -8.8971e-40 + -4.27737e-39 = -5.16708e-39
	(b"00000000011010000101110111001110", b"00000000000000000000000000000000"),
	(b"00000000010010100101110011010101", b"00000000101100101011101010100011"), -- 9.58454e-39 + 6.82913e-39 = 1.64137e-38
	(b"00000000001100000110101110110100", b"00000000000000000000000000000000"),
	(b"00000000001001001111111101001010", b"00000000010101010110101011111110"), -- 4.44674e-39 + 3.39766e-39 = 7.8444e-39
	(b"00000000011001011100010100010001", b"00000000000000000000000000000000"),
	(b"10000000011110110111101101111101", b"10000000000101011011011001101100"), -- 9.34608e-39 + -1.13401e-38 = -1.99399e-39
	(b"00000000001010100111000101001101", b"00000000000000000000000000000000"),
	(b"00000000000011111010011001010010", b"00000000001110100001011110011111"), -- 3.89774e-39 + 1.4372e-39 = 5.33493e-39
	(b"00000000011010000010011001100010", b"00000000000000000000000000000000"),
	(b"10000000011000011101101100011001", b"00000000000001100100101101001001"), -- 9.56466e-39 + -8.98664e-39 = 5.7802e-40
	(b"00000000000011111011101000000011", b"00000000000000000000000000000000"),
	(b"10000000010100010000000110111100", b"10000000010000010100011110111001"), -- 1.44426e-39 + -7.4393e-39 = -5.99504e-39
	(b"00000000000010011101010100111000", b"00000000000000000000000000000000"),
	(b"00000000010000100011110011001100", b"00000000010011000001001000000100"), -- 9.03008e-40 + 6.08295e-39 = 6.98596e-39
	(b"00000000010101000100001001000000", b"00000000000000000000000000000000"),
	(b"10000000000000000110111000111010", b"00000000010100111101010000000110"), -- 7.73795e-39 + -3.95418e-41 = 7.69841e-39
	(b"00000000000100011101111011010101", b"00000000000000000000000000000000"),
	(b"10000000010000110011110101000100", b"10000000001100010101111001101111"), -- 1.64114e-39 + -6.17496e-39 = -4.53382e-39
	(b"00000000010010010010100010000000", b"00000000000000000000000000000000"),
	(b"10000000011001001111011111100001", b"10000000000110111100111101100001"), -- 6.71852e-39 + -9.27247e-39 = -2.55395e-39
	(b"10000000011010111110110111111101", b"00000000000000000000000000000000"),
	(b"10000000001000111100110000001010", b"10000000100011111011101000000111"), -- -9.91177e-39 + -3.28744e-39 = -1.31992e-38
	(b"10000000001100110100101011011101", b"00000000000000000000000000000000"),
	(b"00000000010011100011011000110110", b"00000000000110101110101101011001"), -- -4.71047e-39 + 7.18262e-39 = 2.47215e-39
	(b"10000000001110001101110110001110", b"00000000000000000000000000000000"),
	(b"10000000011000110011001010111101", b"10000000100111000001000001001011"), -- -5.22227e-39 + -9.10992e-39 = -1.43322e-38
	(b"00000000000100001010011001100001", b"00000000000000000000000000000000"),
	(b"10000000010001011011011010010100", b"10000000001101010001000000110011"), -- 1.52905e-39 + -6.40215e-39 = -4.87309e-39
	(b"10000000010010000010101010011000", b"00000000000000000000000000000000"),
	(b"00000000001001010000100101101101", b"10000000001000110010000100101011"), -- -6.62744e-39 + 3.40129e-39 = -3.22614e-39
	(b"00000000001011000010010011111011", b"00000000000000000000000000000000"),
	(b"00000000001100011101010000001000", b"00000000010111011111100100000011"), -- 4.05403e-39 + 4.576e-39 = 8.63003e-39
	(b"10000000000010001011000001010111", b"00000000000000000000000000000000"),
	(b"10000000010100010010110101011000", b"10000000010110011101110110101111"), -- -7.97943e-40 + -7.45494e-39 = -8.25288e-39
	(b"10000000010000001001000010111000", b"00000000000000000000000000000000"),
	(b"10000000010101001011000100101111", b"10000000100101010100000111100111"), -- -5.92939e-39 + -7.77774e-39 = -1.37071e-38
	(b"00000000010110010110110100110000", b"00000000000000000000000000000000"),
	(b"10000000001010001011000111111101", b"00000000001100001011101100110011"), -- 8.21253e-39 + -3.73727e-39 = 4.47526e-39
	(b"00000000010101010001000100110111", b"00000000000000000000000000000000"),
	(b"00000000000100001010011101010000", b"00000000011001011011100010000111"), -- 7.81219e-39 + 1.52939e-39 = 9.34158e-39
	(b"10000000000010111011000010011011", b"00000000000000000000000000000000"),
	(b"10000000001011011000100100011011", b"10000000001110010011100110110110"), -- -1.07354e-39 + -4.18178e-39 = -5.25533e-39
	(b"10000000010111000000110110010110", b"00000000000000000000000000000000"),
	(b"10000000001100001011110000001111", b"10000000100011001100100110100101"), -- -8.45374e-39 + -4.47557e-39 = -1.29293e-38
	(b"10000000001011000001010111000011", b"00000000000000000000000000000000"),
	(b"00000000000010100010010100001001", b"10000000001000011111000010111010"), -- -4.04857e-39 + 9.31641e-40 = -3.11693e-39
	(b"10000000011111000011000010010101", b"00000000000000000000000000000000"),
	(b"00000000010110101001000010011110", b"10000000001000011001111111110111"), -- -1.1405e-38 + 8.31707e-39 = -3.08796e-39
	(b"10000000011010011011000011110000", b"00000000000000000000000000000000"),
	(b"00000000001100110100011011110000", b"10000000001101100110101000000000"), -- -9.7062e-39 + 4.70906e-39 = -4.99714e-39
	(b"10000000011111001100111001110011", b"00000000000000000000000000000000"),
	(b"00000000001000001101010110010011", b"10000000010110111111100011100000"), -- -1.14617e-38 + 3.01535e-39 = -8.44631e-39
	(b"10000000001100011110010111100010", b"00000000000000000000000000000000"),
	(b"10000000000110100111001110111000", b"10000000010011000101100110011010"), -- -4.58241e-39 + -2.42923e-39 = -7.01164e-39
	(b"10000000010111001010101101101111", b"00000000000000000000000000000000"),
	(b"00000000001010111100000010001111", b"10000000001100001110101011100000"), -- -8.51036e-39 + 4.018e-39 = -4.49236e-39
	(b"00000000001011011011000001001111", b"00000000000000000000000000000000"),
	(b"00000000010010101111100101110110", b"00000000011110001010100111000101"), -- 4.19584e-39 + 6.88532e-39 = 1.10812e-38
	(b"10000000001111000101001001110000", b"00000000000000000000000000000000"),
	(b"10000000011001000010110110111010", b"10000000101000001000000000101010"), -- -5.5397e-39 + -9.19995e-39 = -1.47397e-38
	(b"10000000000111110101111101010101", b"00000000000000000000000000000000"),
	(b"10000000001011111001010000111010", b"10000000010011101111001110001111"), -- -2.8811e-39 + -4.36944e-39 = -7.25054e-39
	(b"10000000011110010100000101110101", b"00000000000000000000000000000000"),
	(b"00000000011000111001100110100001", b"10000000000101011010011111010100"), -- -1.11356e-38 + 9.14683e-39 = -1.98875e-39
	(b"10000000001000010001111101001011", b"00000000000000000000000000000000"),
	(b"00000000011100000011101111001111", b"00000000010011110001110010000100"), -- -3.0418e-39 + 1.0307e-38 = 7.26523e-39
	(b"00000000001100000111111101111111", b"00000000000000000000000000000000"),
	(b"00000000011011011101110010101100", b"00000000100111100101110000101011"), -- 4.45384e-39 + 1.00892e-38 = 1.45431e-38
	(b"10000000010001110101011000101000", b"00000000000000000000000000000000"),
	(b"00000000000111101111101000110100", b"10000000001010000101101111110100"), -- -6.55123e-39 + 2.84482e-39 = -3.70641e-39
	(b"00000000011100110001011001001010", b"00000000000000000000000000000000"),
	(b"10000000000011001001100101100110", b"00000000011001100111110011100100"), -- 1.05691e-38 + -1.15705e-39 = 9.41202e-39
	(b"00000000011010100111001010100100", b"00000000000000000000000000000000"),
	(b"10000000010000110111011110000110", b"00000000001001101111101100011110"), -- 9.77569e-39 + -6.19586e-39 = 3.57983e-39
	(b"00000000011000111010100000111100", b"00000000000000000000000000000000"),
	(b"00000000001011111001000001101001", b"00000000100100110011100010100101"), -- 9.15207e-39 + 4.36807e-39 = 1.35201e-38
	(b"10000000011010101000101001000110", b"00000000000000000000000000000000"),
	(b"10000000011100010101100101000100", b"10000000110110111110001110001010"), -- -9.78417e-39 + -1.04094e-38 = -2.01936e-38
	(b"10000000000001100111110110111100", b"00000000000000000000000000000000"),
	(b"10000000001001001010101110100010", b"10000000001010110010100101011110"), -- -5.96118e-40 + -3.36765e-39 = -3.96377e-39
	(b"00000000000111001001100001010001", b"00000000000000000000000000000000"),
	(b"00000000010100010100101111000100", b"00000000011011011110010000010101"), -- 2.62603e-39 + 7.46585e-39 = 1.00919e-38
	(b"00000000010000000100010110011101", b"00000000000000000000000000000000"),
	(b"00000000011110111001111111111010", b"00000000101110111110010110010111"), -- 5.90244e-39 + 1.13532e-38 = 1.72556e-38
	(b"00000000000101011100001011100000", b"00000000000000000000000000000000"),
	(b"00000000011000100110100101010001", b"00000000011110000010110000110001"), -- 1.99845e-39 + 9.03766e-39 = 1.10361e-38
	(b"00000000011111110000010001010110", b"00000000000000000000000000000000"),
	(b"10000000001111110011110001001101", b"00000000001111111100100000001001"), -- 1.16647e-38 + -5.80727e-39 = 5.8574e-39
	(b"10000000011101110010101100110110", b"00000000000000000000000000000000"),
	(b"10000000000011100111110111000001", b"10000000100001011010100011110111"), -- -1.09439e-38 + -1.33081e-39 = -1.22747e-38
	(b"00000000011001001010111010010101", b"00000000000000000000000000000000"),
	(b"00000000000100011001000000111010", b"00000000011101100011111011001111"), -- 9.24618e-39 + 1.61294e-39 = 1.08591e-38
	(b"10000000010111011111100011110111", b"00000000000000000000000000000000"),
	(b"10000000001000011010101000010101", b"10000000011111111010001100001100"), -- -8.63001e-39 + -3.09159e-39 = -1.17216e-38
	(b"00000000011010000010110001000011", b"00000000000000000000000000000000"),
	(b"00000000000010000011010001011000", b"00000000011100000110000010011011"), -- 9.56677e-39 + 7.53461e-40 = 1.03202e-38
	(b"00000000011101100100110101000000", b"00000000000000000000000000000000"),
	(b"00000000001001111001111010100011", b"00000000100111011110101111100011"), -- 1.08643e-38 + 3.63849e-39 = 1.45028e-38
	(b"10000000010101000000001100000010", b"00000000000000000000000000000000"),
	(b"00000000000100011010000000100011", b"10000000010000100110001011011111"), -- -7.71526e-39 + 1.61865e-39 = -6.09661e-39
	(b"00000000010111111101100100110100", b"00000000000000000000000000000000"),
	(b"00000000001011111000011010000110", b"00000000100011110101111110111010"), -- 8.80229e-39 + 4.36453e-39 = 1.31668e-38
	(b"10000000000000001001000101010101", b"00000000000000000000000000000000"),
	(b"00000000010110110110110000101011", b"00000000010110101101101011010110"), -- -5.21353e-41 + 8.39583e-39 = 8.3437e-39
	(b"00000000010101011010100011010011", b"00000000000000000000000000000000"),
	(b"10000000011000110111001111001101", b"10000000000011011100101011111010"), -- 7.86658e-39 + -9.13326e-39 = -1.26668e-39
	(b"00000000000111010011001110000001", b"00000000000000000000000000000000"),
	(b"10000000011100011010101011010000", b"10000000010101000111011101001111"), -- 2.68171e-39 + -1.04387e-38 = -7.75698e-39
	(b"10000000001000010100100000100001", b"00000000000000000000000000000000"),
	(b"00000000000001001010111111101101", b"10000000000111001001100000110100"), -- -3.05645e-39 + 4.30452e-40 = -2.62599e-39
	(b"10000000011000111011110010101001", b"00000000000000000000000000000000"),
	(b"00000000010100111101010011001111", b"10000000000011111110011111011010"), -- -9.15939e-39 + 7.69869e-39 = -1.46071e-39
	(b"00000000000100100011000001110100", b"00000000000000000000000000000000"),
	(b"10000000010111110111011010111000", b"10000000010011010100011001000100"), -- 1.67042e-39 + -8.76696e-39 = -7.09654e-39
	(b"10000000001110111111111110010001", b"00000000000000000000000000000000"),
	(b"00000000000011101101001011010111", b"10000000001011010010110010111010"), -- -5.50997e-39 + 1.36133e-39 = -4.14864e-39
	(b"00000000010100110110001100100010", b"00000000000000000000000000000000"),
	(b"10000000000100010001010110000100", b"00000000010000100100110110011110"), -- 7.65791e-39 + -1.56892e-39 = 6.08899e-39
	(b"00000000011110111100110101011110", b"00000000000000000000000000000000"),
	(b"10000000010000110101001011101100", b"00000000001110000111101001110010"), -- 1.13694e-38 + -6.18273e-39 = 5.18671e-39
	(b"10000000001100110101001011001000", b"00000000000000000000000000000000"),
	(b"00000000000000101001000011001111", b"10000000001100001100000111111001"), -- -4.71331e-39 + 2.35619e-40 = -4.47769e-39
	(b"10000000001100000111011110011001", b"00000000000000000000000000000000"),
	(b"00000000011100011110100001000111", b"00000000010000010111000010101110"), -- -4.45101e-39 + 1.04607e-38 = 6.00973e-39
	(b"00000000011000110110100000011000", b"00000000000000000000000000000000"),
	(b"10000000011010000001010001100011", b"10000000000001001010110001001011"), -- 9.12906e-39 + -9.5582e-39 = -4.29149e-40
	(b"00000000011001111010011111011100", b"00000000000000000000000000000000"),
	(b"00000000010001101011110011101101", b"00000000101011100110010011001001"), -- 9.51927e-39 + 6.49626e-39 = 1.60155e-38
	(b"00000000000101010001001111100011", b"00000000000000000000000000000000"),
	(b"00000000011011000100001000000000", b"00000000100000010101010111100011"), -- 1.93568e-39 + 9.94191e-39 = 1.18776e-38
	(b"10000000001000110010110010000001", b"00000000000000000000000000000000"),
	(b"10000000011010110011111100101000", b"10000000100011100110101110101001"), -- -3.23021e-39 + -9.84905e-39 = -1.30793e-38
	(b"10000000011000011100110110110001", b"00000000000000000000000000000000"),
	(b"10000000010101101111011101001001", b"10000000101110001100010011111010"), -- -8.98183e-39 + -7.98656e-39 = -1.69684e-38
	(b"10000000010100101110001110001111", b"00000000000000000000000000000000"),
	(b"10000000010011100111110011110110", b"10000000101000010110000010000101"), -- -7.61214e-39 + -7.208e-39 = -1.48201e-38
	(b"10000000001110010001010010001011", b"00000000000000000000000000000000"),
	(b"00000000000010010101000011110110", b"10000000001011111100001110010101"), -- -5.24199e-39 + 8.55563e-40 = -4.38643e-39
	(b"10000000001100110100010110001100", b"00000000000000000000000000000000"),
	(b"10000000010100100001101111101100", b"10000000100001010110000101111000"), -- -4.70856e-39 + -7.54053e-39 = -1.22491e-38
	(b"10000000010011101010011000011111", b"00000000000000000000000000000000"),
	(b"10000000001011101000101010101110", b"10000000011111010011000011001101"), -- -7.22276e-39 + -4.27418e-39 = -1.14969e-38
	(b"00000000000101111001111111000100", b"00000000000000000000000000000000"),
	(b"00000000010010000101010001110010", b"00000000010111111111010000110110"), -- 2.16953e-39 + 6.64245e-39 = 8.81198e-39
	(b"00000000000111100011010111000110", b"00000000000000000000000000000000"),
	(b"00000000010000001100011011110100", b"00000000010111101111110010111010"), -- 2.77436e-39 + 5.94884e-39 = 8.7232e-39
	(b"10000000001111111111110110110000", b"00000000000000000000000000000000"),
	(b"10000000010010100011011101011011", b"10000000100010100011010100001011"), -- -5.87664e-39 + -6.81568e-39 = -1.26923e-38
	(b"10000000010101010111110010100001", b"00000000000000000000000000000000"),
	(b"00000000001111000101011011001010", b"10000000000110010010010111010111"), -- -7.85073e-39 + 5.54126e-39 = -2.30946e-39
	(b"10000000010111110101011100111110", b"00000000000000000000000000000000"),
	(b"00000000001101000010011001111111", b"10000000001010110011000010111111"), -- -8.75567e-39 + 4.78926e-39 = -3.96641e-39
	(b"00000000011011011010010100110111", b"00000000000000000000000000000000"),
	(b"00000000000100110100111110110011", b"00000000100000001111010011101010"), -- 1.00693e-38 + 1.77347e-39 = 1.18428e-38
	(b"10000000011001101111100010100010", b"00000000000000000000000000000000"),
	(b"10000000010010101100011110101011", b"10000000101100011100000001001101"), -- -9.45641e-39 + -6.86745e-39 = -1.63239e-38
	(b"00000000010110011100000110010101", b"00000000000000000000000000000000"),
	(b"10000000010001000100110111011011", b"00000000000101010111001110111010"), -- 8.2428e-39 + -6.27274e-39 = 1.97006e-39
	(b"10000000000010010111110100101011", b"00000000000000000000000000000000"),
	(b"10000000000010000111001000000100", b"10000000000100011110111100101111"), -- -8.71421e-40 + -7.75585e-40 = -1.64701e-39
	(b"00000000001110110100101101001110", b"00000000000000000000000000000000"),
	(b"00000000001111110010111101100001", b"00000000011110100111101010101111"), -- 5.44531e-39 + 5.80263e-39 = 1.12479e-38
	(b"10000000010000101001001100110000", b"00000000000000000000000000000000"),
	(b"10000000011101110011100001010111", b"10000000101110011100101110000111"), -- -6.11394e-39 + -1.09486e-38 = -1.70626e-38
	(b"10000000001100011011001110111101", b"00000000000000000000000000000000"),
	(b"00000000001110000101111000111101", b"00000000000001101010101010000000"), -- -4.56442e-39 + 5.17659e-39 = 6.12177e-40
	(b"10000000001010111010110011101110", b"00000000000000000000000000000000"),
	(b"00000000010001100000000110110010", b"00000000000110100101010011000100"), -- -4.01096e-39 + 6.42909e-39 = 2.41813e-39
	(b"00000000011001100001000101000000", b"00000000000000000000000000000000"),
	(b"00000000001111100101110000101000", b"00000000101001000110110101101000"), -- 9.37341e-39 + 5.72686e-39 = 1.51003e-38
	(b"10000000011001000010001101001110", b"00000000000000000000000000000000"),
	(b"10000000000111010110000010000101", b"10000000100000011000001111010011"), -- -9.19621e-39 + -2.69785e-39 = -1.18941e-38
	(b"10000000010010001101011110011101", b"00000000000000000000000000000000"),
	(b"00000000001001110010110010110010", b"10000000001000011010101011101011"), -- -6.6895e-39 + 3.59762e-39 = -3.09189e-39
	(b"10000000010001011101011110101001", b"00000000000000000000000000000000"),
	(b"00000000010100101101001000101001", b"00000000000011001111101010000000"), -- -6.41401e-39 + 7.6059e-39 = 1.19189e-39
	(b"00000000001000001011100101100100", b"00000000000000000000000000000000"),
	(b"10000000001111100010100011110010", b"10000000000111010110111110001110"), -- 3.00524e-39 + -5.70849e-39 = -2.70325e-39
	(b"00000000000111010000110010110000", b"00000000000000000000000000000000"),
	(b"00000000010101101001001110000000", b"00000000011100111010000000110000"), -- 2.66778e-39 + 7.95077e-39 = 1.06185e-38
	(b"10000000011010101101011010011100", b"00000000000000000000000000000000"),
	(b"10000000000101010100001011011001", b"10000000100000000001100101110101"), -- -9.81155e-39 + -1.95253e-39 = -1.17641e-38
	(b"00000000011110111011001010111111", b"00000000000000000000000000000000"),
	(b"10000000001110001000000101101010", b"00000000010000110011000101010101"), -- 1.13599e-38 + -5.18921e-39 = 6.17068e-39
	(b"00000000011110011111111011010111", b"00000000000000000000000000000000"),
	(b"10000000010111100110010100111100", b"00000000000110111001100110011011"), -- 1.12035e-38 + -8.66885e-39 = 2.53466e-39
	(b"10000000001111001010011100100110", b"00000000000000000000000000000000"),
	(b"00000000010110100010110100100011", b"00000000000111011000010111111101"), -- -5.57009e-39 + 8.28139e-39 = 2.7113e-39
	(b"10000000010110010111101001111001", b"00000000000000000000000000000000"),
	(b"00000000010000001011110100011111", b"10000000000110001011110101011010"), -- -8.21729e-39 + 5.94532e-39 = -2.27198e-39
	(b"00000000011101001000000000100000", b"00000000000000000000000000000000"),
	(b"10000000000011100000101000100001", b"00000000011001100111010111111111"), -- 1.06989e-38 + -1.28933e-39 = 9.40955e-39
	(b"00000000000100011101011101100010", b"00000000000000000000000000000000"),
	(b"10000000010100111100111010111001", b"10000000010000011111011101010111"), -- 1.63847e-39 + -7.6965e-39 = -6.05804e-39
	(b"10000000000011111001000001000111", b"00000000000000000000000000000000"),
	(b"00000000001110110001010000100111", b"00000000001010111000001111100000"), -- -1.42929e-39 + 5.42552e-39 = 3.99623e-39
	(b"00000000010101000000110110100001", b"00000000000000000000000000000000"),
	(b"00000000010010111010001110000100", b"00000000100111111011000100100101"), -- 7.71907e-39 + 6.94632e-39 = 1.46654e-38
	(b"00000000000000100011100110110010", b"00000000000000000000000000000000"),
	(b"00000000001100111111110011001111", b"00000000001101100011011010000001"), -- 2.04368e-40 + 4.7743e-39 = 4.97867e-39
	(b"00000000011101110100110011111011", b"00000000000000000000000000000000"),
	(b"00000000011100001101100010111110", b"00000000111010000010010110111001"), -- 1.0956e-38 + 1.03633e-38 = 2.13194e-38
	(b"10000000011100110101100101101011", b"00000000000000000000000000000000"),
	(b"10000000000110100001001010011101", b"10000000100011010110110000001000"), -- -1.05932e-38 + -2.3944e-39 = -1.29876e-38
	(b"10000000010100111010011000101011", b"00000000000000000000000000000000"),
	(b"10000000011001111001111011001011", b"10000000101110110100010011110110"), -- -7.68196e-39 + -9.51602e-39 = -1.7198e-38
	(b"00000000001010110110110110101011", b"00000000000000000000000000000000"),
	(b"00000000010111110010111110010001", b"00000000100010101001110100111100"), -- 3.98827e-39 + 8.74144e-39 = 1.27297e-38
	(b"00000000010000111001011101010101", b"00000000000000000000000000000000"),
	(b"10000000011011110111111010110010", b"10000000001010111110011101011101"), -- 6.20727e-39 + -1.02392e-38 = -4.03192e-39
	(b"00000000011111101010011111000111", b"00000000000000000000000000000000"),
	(b"10000000001011111101111011001000", b"00000000010011101100100011111111"), -- 1.16315e-38 + -4.39619e-39 = 7.23527e-39
	(b"00000000000101100111111000011010", b"00000000000000000000000000000000"),
	(b"10000000001101111011111001011001", b"10000000001000010100000000111111"), -- 2.06562e-39 + -5.11924e-39 = -3.05362e-39
	(b"00000000011101110100011011011101", b"00000000000000000000000000000000"),
	(b"00000000001000010001110001100110", b"00000000100110000110001101000011"), -- 1.09538e-38 + 3.04076e-39 = 1.39946e-38
	(b"00000000011000111001101011111001", b"00000000000000000000000000000000"),
	(b"10000000001010101011000010000110", b"00000000001110001110101001110011"), -- 9.14731e-39 + -3.92042e-39 = 5.22689e-39
	(b"00000000000000110101001011101010", b"00000000000000000000000000000000"),
	(b"00000000011000101000111110010100", b"00000000011001011110001001111110"), -- 3.0525e-40 + 9.05138e-39 = 9.35664e-39
	(b"10000000011100111110100010100000", b"00000000000000000000000000000000"),
	(b"00000000011000101010101101101100", b"10000000000100010011110100110100"), -- -1.06445e-38 + 9.06137e-39 = -1.58316e-39
	(b"10000000000101010111001010101101", b"00000000000000000000000000000000"),
	(b"10000000001000110000011010011010", b"10000000001110000111100101000111"), -- -1.96968e-39 + -3.21661e-39 = -5.18629e-39
	(b"00000000010110000110010000101001", b"00000000000000000000000000000000"),
	(b"00000000001000000001101111110010", b"00000000011110001000000000011011"), -- 8.11745e-39 + 2.94876e-39 = 1.10662e-38
	(b"10000000011110101010110110111010", b"00000000000000000000000000000000"),
	(b"10000000001100110001110100011110", b"10000000101011011100101011011000"), -- -1.12663e-38 + -4.69406e-39 = -1.59603e-38
	(b"10000000000001011100000001000110", b"00000000000000000000000000000000"),
	(b"10000000001100010010010101010010", b"10000000001101101110010110011000"), -- -5.28152e-40 + -4.51333e-39 = -5.04148e-39
	(b"10000000011111110100111011101100", b"00000000000000000000000000000000"),
	(b"10000000001110110110010011100000", b"10000000101110101011001111001100"), -- -1.16914e-38 + -5.45448e-39 = -1.71459e-38
	(b"10000000000111100010000110001011", b"00000000000000000000000000000000"),
	(b"00000000010011001001100110010010", b"00000000001011100111100000000111"), -- -2.7671e-39 + 7.03459e-39 = 4.26749e-39
	(b"00000000010111000011001101100101", b"00000000000000000000000000000000"),
	(b"10000000011001011110001010100000", b"10000000000010011010111100111011"), -- 8.4673e-39 + -9.35668e-39 = -8.8938e-40
	(b"10000000000000011010110101001000", b"00000000000000000000000000000000"),
	(b"00000000000110000110011110000011", b"00000000000101101011101000111011"), -- -1.53997e-40 + 2.24118e-39 = 2.08719e-39
	(b"10000000000110100111101000110010", b"00000000000000000000000000000000"),
	(b"10000000011011000110100001000101", b"10000000100001101110001001110111"), -- -2.43156e-39 + -9.95564e-39 = -1.23872e-38
	(b"00000000011000000010010101000100", b"00000000000000000000000000000000"),
	(b"10000000011100000011011100101100", b"10000000000100000001000111101000"), -- 8.82958e-39 + -1.03054e-38 = -1.47579e-39
	(b"00000000001100001101010111001101", b"00000000000000000000000000000000"),
	(b"10000000001001001111011101100110", b"00000000000010111101111001100111"), -- 4.4848e-39 + -3.39483e-39 = 1.08997e-39
	(b"10000000001010110110010011001111", b"00000000000000000000000000000000"),
	(b"10000000001101010111110101100000", b"10000000011000001110001000101111"), -- -3.98509e-39 + -4.91226e-39 = -8.89735e-39
	(b"10000000010010100100000100100011", b"00000000000000000000000000000000"),
	(b"10000000010001000111100110000011", b"10000000100011101011101010100110"), -- -6.81919e-39 + -6.2884e-39 = -1.31076e-38
	(b"10000000011110110011011101111100", b"00000000000000000000000000000000"),
	(b"00000000010010011111111010110001", b"10000000001100010011100011001011"), -- -1.13157e-38 + 6.79536e-39 = -4.52031e-39
	(b"10000000000000011011101111001001", b"00000000000000000000000000000000"),
	(b"00000000001100001111001001001000", b"00000000001011110011011001111111"), -- -1.592e-40 + 4.49502e-39 = 4.33582e-39
	(b"00000000010001110110010101101100", b"00000000000000000000000000000000"),
	(b"10000000000001010011010100011100", b"00000000010000100011000001010000"), -- 6.5567e-39 + -4.7823e-40 = 6.07847e-39
	(b"10000000000111001001101100000011", b"00000000000000000000000000000000"),
	(b"00000000000101011001101001000111", b"10000000000001110000000010111100"), -- -2.627e-39 + 1.98389e-39 = -6.43112e-40
	(b"00000000011010000001100010000111", b"00000000000000000000000000000000"),
	(b"00000000000101111011010110001110", b"00000000011111111100111000010101"), -- 9.55969e-39 + 2.17735e-39 = 1.1737e-38
	(b"00000000010100111101000000011110", b"00000000000000000000000000000000"),
	(b"10000000000011000101010110001111", b"00000000010001110111101010001111"), -- 7.697e-39 + -1.13272e-39 = 6.56429e-39
	(b"00000000010111001110111100100100", b"00000000000000000000000000000000"),
	(b"00000000010001010110110101100100", b"00000000101000100101110010001000"), -- 8.53465e-39 + 6.37589e-39 = 1.49105e-38
	(b"00000000001111000011101011110010", b"00000000000000000000000000000000"),
	(b"00000000011101111010011011100100", b"00000000101100111110000111010110"), -- 5.53128e-39 + 1.09883e-38 = 1.65196e-38
	(b"10000000011111001101101011001111", b"00000000000000000000000000000000"),
	(b"00000000000110011100111111000000", b"10000000011000110000101100001111"), -- -1.14661e-38 + 2.37041e-39 = -9.09568e-39
	(b"00000000000001010010111010101010", b"00000000000000000000000000000000"),
	(b"00000000011101100001110100001001", b"00000000011110110100101110110011"), -- 4.75917e-40 + 1.0847e-38 = 1.13229e-38
	(b"10000000010000010110101010010100", b"00000000000000000000000000000000"),
	(b"10000000011100010111110111011100", b"10000000101100101110100001110000"), -- -6.00754e-39 + -1.04226e-38 = -1.64301e-38
	(b"10000000001000011110001011101110", b"00000000000000000000000000000000"),
	(b"10000000010001010111100000111001", b"10000000011001110101101100100111"), -- -3.11198e-39 + -6.37978e-39 = -9.49176e-39
	(b"10000000001001111111001001110010", b"00000000000000000000000000000000"),
	(b"00000000010110100010101101111100", b"00000000001100100011100100001010"), -- -3.66856e-39 + 8.28079e-39 = 4.61224e-39
	(b"10000000000111000010111010001010", b"00000000000000000000000000000000"),
	(b"00000000000011110000100101000011", b"10000000000011010010010101000111"), -- -2.58809e-39 + 1.38085e-39 = -1.20723e-39
	(b"00000000010110011100001110010111", b"00000000000000000000000000000000"),
	(b"00000000001111101011110000101101", b"00000000100110000111111111000100"), -- 8.24352e-39 + 5.76131e-39 = 1.40048e-38
	(b"00000000000010000000000101100110", b"00000000000000000000000000000000"),
	(b"00000000000001001110101001111100", b"00000000000011001110101111100010"), -- 7.35186e-40 + 4.51459e-40 = 1.18664e-39
	(b"00000000001011010010001011101101", b"00000000000000000000000000000000"),
	(b"00000000010111111010100010110110", b"00000000100011001100101110100011"), -- 4.14513e-39 + 8.78489e-39 = 1.293e-38
	(b"10000000001111111011111011101001", b"00000000000000000000000000000000"),
	(b"00000000010100111100100001011100", b"00000000000101000000100101110011"), -- -5.85412e-39 + 7.69422e-39 = 1.8401e-39
	(b"00000000010111000110000110100000", b"00000000000000000000000000000000"),
	(b"10000000001011010000101100100011", b"00000000001011110101011001111101"), -- 8.48389e-39 + -4.13659e-39 = 4.34729e-39
	(b"00000000000101010000011101111101", b"00000000000000000000000000000000"),
	(b"00000000000001110000000000010000", b"00000000000111000000011110001101"), -- 1.93123e-39 + 6.42871e-40 = 2.5741e-39
	(b"10000000011001100001101010000111", b"00000000000000000000000000000000"),
	(b"00000000010110000011110011000000", b"10000000000011011101110111000111"), -- -9.37674e-39 + 8.10332e-39 = -1.27342e-39
	(b"10000000011110011101011101101101", b"00000000000000000000000000000000"),
	(b"00000000010000010010010001011100", b"10000000001110001011001100010001"), -- -1.11894e-38 + 5.98235e-39 = -5.20702e-39
	(b"00000000011001010001100000000001", b"00000000000000000000000000000000"),
	(b"10000000011111111111101011011001", b"10000000000110101110001011011000"), -- 9.284e-39 + -1.17531e-38 = -2.4691e-39
	(b"10000000010010000111000000001110", b"00000000000000000000000000000000"),
	(b"10000000010110010110000110011011", b"10000000101000011101000110101001"), -- -6.65235e-39 + -8.20837e-39 = -1.48607e-38
	(b"10000000011110001011001010101110", b"00000000000000000000000000000000"),
	(b"10000000011101100101110111010011", b"10000000111011110001000010000001"), -- -1.10844e-38 + -1.08702e-38 = -2.19546e-38
	(b"10000000000110001100110101010111", b"00000000000000000000000000000000"),
	(b"00000000000110110010101000000001", b"00000000000000100101110010101010"), -- -2.27771e-39 + 2.49463e-39 = 2.16913e-40
	(b"10000000010001110011011110011110", b"00000000000000000000000000000000"),
	(b"00000000010111011011110011110101", b"00000000000101101000010101010111"), -- -6.54027e-39 + 8.60849e-39 = 2.06821e-39
	(b"00000000001101110000001110011001", b"00000000000000000000000000000000"),
	(b"10000000011100100011111100011100", b"10000000001110110011101110000011"), -- 5.05224e-39 + -1.04919e-38 = -5.43964e-39
	(b"00000000000101001010001100101001", b"00000000000000000000000000000000"),
	(b"10000000001111001100011111011011", b"10000000001010000010010010110010"), -- 1.89524e-39 + -5.58182e-39 = -3.68658e-39
	(b"10000000011100000011110111111000", b"00000000000000000000000000000000"),
	(b"10000000001001111111101101111001", b"10000000100110000011100101110001"), -- -1.03078e-38 + -3.6718e-39 = -1.39796e-38
	(b"10000000011010011000111010100110", b"00000000000000000000000000000000"),
	(b"00000000010011001001110111111010", b"10000000000111001111000010101100"), -- -9.6939e-39 + 7.03617e-39 = -2.65773e-39
	(b"00000000001000100001101100110001", b"00000000000000000000000000000000"),
	(b"00000000010011100111001001111011", b"00000000011100001000110110101100"), -- 3.13216e-39 + 7.20424e-39 = 1.03364e-38
	(b"10000000011100110001110001111001", b"00000000000000000000000000000000"),
	(b"00000000001001101101110110111111", b"10000000010011000011111010111010"), -- -1.05713e-38 + 3.5693e-39 = -7.002e-39
	(b"00000000001110001110010010011101", b"00000000000000000000000000000000"),
	(b"10000000001001000110100111100011", b"00000000000101000111101010111010"), -- 5.2248e-39 + -3.34406e-39 = 1.88074e-39
	(b"00000000000001010010110011110010", b"00000000000000000000000000000000"),
	(b"10000000001001111010110011011010", b"10000000001000100111111111101000"), -- 4.75301e-40 + -3.64359e-39 = -3.16829e-39
	(b"10000000010101000100100010010000", b"00000000000000000000000000000000"),
	(b"00000000010111001000101000010110", b"00000000000010000100000110000110"), -- -7.74021e-39 + 8.4984e-39 = 7.58189e-40
	(b"00000000001010000111110010001011", b"00000000000000000000000000000000"),
	(b"00000000011011111110000000001111", b"00000000100110000101110010011010"), -- 3.7181e-39 + 1.02741e-38 = 1.39922e-38
	(b"00000000001011011100010000011110", b"00000000000000000000000000000000"),
	(b"10000000000011110111110010110111", b"00000000000111100100011101100111"), -- 4.20295e-39 + -1.42227e-39 = 2.78068e-39
	(b"10000000001001010110101111010101", b"00000000000000000000000000000000"),
	(b"10000000010000000001010001110001", b"10000000011001011000000001000110"), -- -3.4366e-39 + -5.8848e-39 = -9.3214e-39
	(b"00000000011010010111110111001011", b"00000000000000000000000000000000"),
	(b"00000000010010111101010001101111", b"00000000101101010101001000111010"), -- 9.68785e-39 + 6.96387e-39 = 1.66517e-38
	(b"00000000011010011100000100010001", b"00000000000000000000000000000000"),
	(b"10000000000011010000110100100000", b"00000000010111001011001111110001"), -- 9.71199e-39 + -1.19857e-39 = 8.51342e-39
	(b"10000000011101001101110100011111", b"00000000000000000000000000000000"),
	(b"10000000010111000000110110011001", b"10000000110100001110101010111000"), -- -1.07322e-38 + -8.45374e-39 = -1.9186e-38
	(b"00000000001111011111001000010010", b"00000000000000000000000000000000"),
	(b"00000000000011110100000001110110", b"00000000010011010011001010001000"), -- 5.6888e-39 + 1.40066e-39 = 7.08946e-39
	(b"10000000010100011111111111001111", b"00000000000000000000000000000000"),
	(b"00000000011000010101110010110101", b"00000000000011110101110011100110"), -- -7.53044e-39 + 8.9413e-39 = 1.41086e-39
	(b"10000000000001100110111011100111", b"00000000000000000000000000000000"),
	(b"00000000011001111110010010000111", b"00000000011000010111010110100000"), -- -5.90797e-40 + 9.54104e-39 = 8.95024e-39
	(b"10000000011100000111010011010110", b"00000000000000000000000000000000"),
	(b"00000000001011011101000011111000", b"10000000010000101010001111011110"), -- -1.03275e-38 + 4.20756e-39 = -6.11993e-39
	(b"10000000011101101000110010100011", b"00000000000000000000000000000000"),
	(b"00000000011001110010101100110010", b"10000000000011110110000101110001"), -- -1.0887e-38 + 9.47455e-39 = -1.41249e-39
	(b"10000000001110110110101111110001", b"00000000000000000000000000000000"),
	(b"00000000000001011010000111011110", b"10000000001101011100101000010011"), -- -5.45702e-39 + 5.17244e-40 = -4.93977e-39
	(b"10000000001001010110111110000111", b"00000000000000000000000000000000"),
	(b"00000000011100110111110000101011", b"00000000010011100000110010100100"), -- -3.43792e-39 + 1.06056e-38 = 7.1677e-39
	(b"00000000000001110100010111111100", b"00000000000000000000000000000000"),
	(b"10000000000100101111101000110110", b"10000000000010111011010000111010"), -- 6.67954e-40 + -1.7428e-39 = -1.07484e-39
	(b"00000000011111000100000111110100", b"00000000000000000000000000000000"),
	(b"10000000000010111011000111111100", b"00000000011100001000111111111000"), -- 1.14113e-38 + -1.07404e-39 = 1.03372e-38
	(b"10000000001101010001001011110010", b"00000000000000000000000000000000"),
	(b"00000000000110011010101111110010", b"10000000000110110110011100000000"), -- -4.87408e-39 + 2.35757e-39 = -2.51651e-39
	(b"10000000000000011000001100101000", b"00000000000000000000000000000000"),
	(b"10000000010011010100101001110100", b"10000000010011101100110110011100"), -- -1.38885e-40 + -7.09804e-39 = -7.23693e-39
	(b"10000000011111001001000000011010", b"00000000000000000000000000000000"),
	(b"10000000010010110110111010101001", b"10000000110001111111111011000011"), -- -1.14393e-38 + -6.92736e-39 = -1.83667e-38
	(b"00000000010110011101111010001110", b"00000000000000000000000000000000"),
	(b"10000000000111010111101111010011", b"00000000001111000110001010111011"), -- 8.2532e-39 + -2.70765e-39 = 5.54555e-39
	(b"10000000010011011011011100100111", b"00000000000000000000000000000000"),
	(b"00000000001000000011100110001110", b"10000000001011010111110110011001"), -- -7.13704e-39 + 2.95938e-39 = -4.17765e-39
	(b"00000000011101100011111010011001", b"00000000000000000000000000000000"),
	(b"00000000000010000111001000110011", b"00000000011111101011000011001100"), -- 1.0859e-38 + 7.75651e-40 = 1.16347e-38
	(b"10000000011000101011111000100110", b"00000000000000000000000000000000"),
	(b"00000000000101011010001101101100", b"10000000010011010001101010111010"), -- -9.06809e-39 + 1.98717e-39 = -7.08092e-39
	(b"00000000001101011001110110100001", b"00000000000000000000000000000000"),
	(b"10000000001010100110100001000000", b"00000000000010110011010101100001"), -- 4.92383e-39 + -3.89449e-39 = 1.02934e-39
	(b"10000000000001000011011111101100", b"00000000000000000000000000000000"),
	(b"00000000011000101101001111110111", b"00000000010111101001110000001011"), -- -3.87403e-40 + 9.07592e-39 = 8.68851e-39
	(b"00000000001111110100100001110011", b"00000000000000000000000000000000"),
	(b"10000000001111001000101100001110", b"00000000000000101011110101100101"), -- 5.81163e-39 + -5.56001e-39 = 2.51613e-40
	(b"10000000010111011110101100000101", b"00000000000000000000000000000000"),
	(b"10000000011110101001011101110111", b"10000000110110001000001001111100"), -- -8.62501e-39 + -1.12583e-38 = -1.98833e-38
	(b"10000000000111011001101010001111", b"00000000000000000000000000000000"),
	(b"10000000010110010000011001010101", b"10000000011101101010000011100100"), -- -2.71867e-39 + -8.17563e-39 = -1.08943e-38
	(b"10000000011000000001110000101101", b"00000000000000000000000000000000"),
	(b"00000000010011101010011000001010", b"10000000000100010111011000100011"), -- -8.82632e-39 + 7.22273e-39 = -1.60358e-39
	(b"10000000000101000100010110101001", b"00000000000000000000000000000000"),
	(b"10000000011001001000101111100010", b"10000000011110001101000110001011"), -- -1.8617e-39 + -9.23373e-39 = -1.10954e-38
	(b"00000000011101010110111101000101", b"00000000000000000000000000000000"),
	(b"00000000000011100111011000010110", b"00000000100000111110010101011011"), -- 1.07847e-38 + 1.32806e-39 = 1.21127e-38
	(b"10000000011010110110011010110110", b"00000000000000000000000000000000"),
	(b"00000000000101011011010011010001", b"10000000010101011011000111100101"), -- -9.86324e-39 + 1.99341e-39 = -7.86983e-39
	(b"10000000001010010001111111101000", b"00000000000000000000000000000000"),
	(b"10000000001011101011000000010010", b"10000000010101111100111111111010"), -- -3.7767e-39 + -4.28759e-39 = -8.0643e-39
	(b"10000000010100000100000100000001", b"00000000000000000000000000000000"),
	(b"00000000010111000001011111000011", b"00000000000010111101011011000010"), -- -7.37016e-39 + 8.45739e-39 = 1.08723e-39
	(b"00000000001101010010000010000010", b"00000000000000000000000000000000"),
	(b"00000000000010001011100010011011", b"00000000001111011101100100011101"), -- 4.87894e-39 + 8.00908e-40 = 5.67985e-39
	(b"10000000000100001000100000110000", b"00000000000000000000000000000000"),
	(b"00000000001111010110110110101010", b"00000000001011001110010101111010"), -- -1.51822e-39 + 5.64131e-39 = 4.12308e-39
	(b"10000000000011000101111010000010", b"00000000000000000000000000000000"),
	(b"10000000001100001100010010110101", b"10000000001111010010001100110111"), -- -1.13593e-39 + -4.47867e-39 = -5.6146e-39
	(b"10000000010001100011000001100100", b"00000000000000000000000000000000"),
	(b"00000000000110010011100001100111", b"10000000001011001111011111111101"), -- -6.44584e-39 + 2.31612e-39 = -4.12972e-39
	(b"10000000000111101010110110000001", b"00000000000000000000000000000000"),
	(b"10000000000100100010001000111110", b"10000000001100001100111110111111"), -- -2.81731e-39 + -1.66532e-39 = -4.48263e-39
	(b"10000000011100000010000101011100", b"00000000000000000000000000000000"),
	(b"00000000011101010101100010000011", b"00000000000001010011011100100111"), -- -1.02975e-38 + 1.07765e-38 = 4.78962e-40
	(b"00000000000000101100011111101001", b"00000000000000000000000000000000"),
	(b"00000000011010111001100110011110", b"00000000011011100110000110000111"), -- 2.55385e-40 + 9.88151e-39 = 1.01369e-38
	(b"00000000000110101110010101010010", b"00000000000000000000000000000000"),
	(b"10000000011100011001010100110011", b"10000000010101101010111111100001"), -- 2.46999e-39 + -1.04309e-38 = -7.96095e-39
	(b"00000000010011110110101011111110", b"00000000000000000000000000000000"),
	(b"10000000011111100011011000101011", b"10000000001011101100101100101101"), -- 7.29339e-39 + -1.15907e-38 = -4.29732e-39
	(b"00000000000011111110001001110000", b"00000000000000000000000000000000"),
	(b"10000000011111010110101000001111", b"10000000011011011000011110011111"), -- 1.45876e-39 + -1.15175e-38 = -1.00587e-38
	(b"00000000000110001010110110010001", b"00000000000000000000000000000000"),
	(b"00000000001100001011001010110111", b"00000000010010010110000001001000"), -- 2.26632e-39 + 4.47221e-39 = 6.73853e-39
	(b"10000000000100110111101101010001", b"00000000000000000000000000000000"),
	(b"00000000000111011101010001001010", b"00000000000010100101100011111001"), -- -1.78911e-39 + 2.73938e-39 = 9.50272e-40
	(b"10000000000111111111100010110110", b"00000000000000000000000000000000"),
	(b"10000000011111111001111101000011", b"10000000100111111001011111111001"), -- -2.93612e-39 + -1.17202e-38 = -1.46564e-38
	(b"00000000001110010111011000100010", b"00000000000000000000000000000000"),
	(b"10000000001100101001100010101011", b"00000000000001101101110101110111"), -- 5.277e-39 + -4.64654e-39 = 6.3046e-40
	(b"00000000000001000011011000111111", b"00000000000000000000000000000000"),
	(b"00000000001000010011100110101010", b"00000000001001010110111111101001"), -- 3.86802e-40 + 3.05126e-39 = 3.43806e-39
	(b"00000000000101100100111111000111", b"00000000000000000000000000000000"),
	(b"10000000001111010011100000000101", b"10000000001001101110100000111110"), -- 2.049e-39 + -5.62206e-39 = -3.57306e-39
	(b"00000000001110010110010111110100", b"00000000000000000000000000000000"),
	(b"10000000010001100010001100111011", b"10000000000011001011110101000111"), -- 5.2712e-39 + -6.44112e-39 = -1.16993e-39
	(b"10000000010010001011001111001100", b"00000000000000000000000000000000"),
	(b"00000000001100101000000111110010", b"10000000000101100011000111011010"), -- -6.67665e-39 + 4.63839e-39 = -2.03826e-39
	(b"00000000001110100110101100111111", b"00000000000000000000000000000000"),
	(b"10000000010000000110111100100110", b"10000000000001100000001111100111"), -- 5.36493e-39 + -5.91734e-39 = -5.52413e-40
	(b"00000000011000010111000110101001", b"00000000000000000000000000000000"),
	(b"10000000001100111101010110011101", b"00000000001011011001110000001100"), -- 8.94882e-39 + -4.76024e-39 = 4.18858e-39
	(b"10000000000011010101111000001111", b"00000000000000000000000000000000"),
	(b"10000000000100000111101000010100", b"10000000000111011101100000100011"), -- -1.2276e-39 + -1.51316e-39 = -2.74076e-39
	(b"10000000011110100100111000111001", b"00000000000000000000000000000000"),
	(b"00000000011010000111100010001110", b"10000000000100011101010110101011"), -- -1.1232e-38 + 9.59414e-39 = -1.63785e-39
	(b"10000000011100011001111011011111", b"00000000000000000000000000000000"),
	(b"00000000010111110011100000001100", b"10000000000100100110011011010011"), -- -1.04344e-38 + 8.74448e-39 = -1.68993e-39
	(b"00000000011100001011010000110010", b"00000000000000000000000000000000"),
	(b"10000000010011001101011110010111", b"00000000001000111101110010011011"), -- 1.03502e-38 + -7.05684e-39 = 3.29338e-39
	(b"00000000011001110001101001011000", b"00000000000000000000000000000000"),
	(b"00000000001000000000101010010001", b"00000000100001110010010011101001"), -- 9.46851e-39 + 2.94253e-39 = 1.2411e-38
	(b"10000000000110001100011101101001", b"00000000000000000000000000000000"),
	(b"10000000000100110110100011000011", b"10000000001011000011000000101100"), -- -2.27559e-39 + -1.78246e-39 = -4.05804e-39
	(b"10000000000010110111110001000101", b"00000000000000000000000000000000"),
	(b"10000000011101111101111011000010", b"10000000100000110101101100000111"), -- -1.05477e-39 + -1.10083e-38 = -1.20631e-38
	(b"10000000000100001100001100011101", b"00000000000000000000000000000000"),
	(b"00000000010111000100101011100010", b"00000000010010111000011111000101"), -- -1.53936e-39 + 8.47573e-39 = 6.93637e-39
	(b"10000000010000001101011111101110", b"00000000000000000000000000000000"),
	(b"00000000001011100101010101010110", b"10000000000100101000001010011000"), -- -5.95493e-39 + 4.25505e-39 = -1.69989e-39
	(b"00000000001111100000001110011011", b"00000000000000000000000000000000"),
	(b"10000000000101010110001101001010", b"00000000001010001010000001010001"), -- 5.69509e-39 + -1.96416e-39 = 3.73093e-39
	(b"00000000000001100110111001010001", b"00000000000000000000000000000000"),
	(b"10000000000011010010001101101100", b"10000000000001101011010100011011"), -- 5.90587e-40 + -1.20657e-39 = -6.15981e-40
	(b"10000000001000010000010011011011", b"00000000000000000000000000000000"),
	(b"10000000010000100010101010110000", b"10000000011000110010111110001011"), -- -3.03231e-39 + -6.07646e-39 = -9.10877e-39
	(b"10000000000100010111111101111000", b"00000000000000000000000000000000"),
	(b"10000000010111011011101001110000", b"10000000011011110011100111101000"), -- -1.60693e-39 + -8.60758e-39 = -1.02145e-38
	(b"00000000011000000010001100100111", b"00000000000000000000000000000000"),
	(b"00000000011101001111011000000111", b"00000000110101010001100100101110"), -- 8.82882e-39 + 1.07412e-38 = 1.957e-38
	(b"00000000000111111000001110011101", b"00000000000000000000000000000000"),
	(b"00000000000101000001101001101100", b"00000000001100111001111000001001"), -- 2.89411e-39 + 1.84619e-39 = 4.7403e-39
	(b"00000000001101011101001110101111", b"00000000000000000000000000000000"),
	(b"00000000001110000011101010000010", b"00000000011011100000111000110001"), -- 4.94322e-39 + 5.16378e-39 = 1.0107e-38
	(b"00000000000111011100010010101110", b"00000000000000000000000000000000"),
	(b"10000000010010010010010101100110", b"10000000001010110110000010111000"), -- 2.73378e-39 + -6.71741e-39 = -3.98362e-39
	(b"10000000010111000010000101010010", b"00000000000000000000000000000000"),
	(b"00000000001000001000000001110001", b"10000000001110111010000011100001"), -- -8.46082e-39 + 2.98481e-39 = -5.47601e-39
	(b"10000000000011111101000101100101", b"00000000000000000000000000000000"),
	(b"00000000010110101001110111000010", b"00000000010010101100110001011101"), -- -1.45265e-39 + 8.32179e-39 = 6.86914e-39
	(b"10000000001110101110110101111101", b"00000000000000000000000000000000"),
	(b"10000000010011110110101110001110", b"10000000100010100101100100001011"), -- -5.41165e-39 + -7.29359e-39 = -1.27052e-38
	(b"00000000010111100010100001011111", b"00000000000000000000000000000000"),
	(b"10000000001010010101110001010011", b"00000000001101001100110000001100"), -- 8.64702e-39 + -3.79838e-39 = 4.84864e-39
	(b"10000000000000101101100010101111", b"00000000000000000000000000000000"),
	(b"00000000010011011100011100010011", b"00000000010010101110111001100100"), -- -2.61402e-40 + 7.14275e-39 = 6.88135e-39
	(b"00000000010010110111011111101000", b"00000000000000000000000000000000"),
	(b"00000000011111011010111101101101", b"00000000110010010010011101010101"), -- 6.93068e-39 + 1.15424e-38 = 1.8473e-38
	(b"10000000000011110001001011011001", b"00000000000000000000000000000000"),
	(b"00000000001011111100101011101111", b"00000000001000001011100000010110"), -- -1.38429e-39 + 4.38907e-39 = 3.00477e-39
	(b"00000000000110110110011111001010", b"00000000000000000000000000000000"),
	(b"10000000000100111110000101111011", b"00000000000001111000011001001111"), -- 2.51679e-39 + -1.82576e-39 = 6.91029e-40
	(b"10000000001101001111000000011001", b"00000000000000000000000000000000"),
	(b"10000000001100001011100001000001", b"10000000011001011010100001011010"), -- -4.86158e-39 + -4.4742e-39 = -9.33578e-39
	(b"00000000010011100011111001111110", b"00000000000000000000000000000000"),
	(b"00000000000001100001000000010110", b"00000000010101000100111010010100"), -- 7.18559e-39 + 5.56784e-40 = 7.74237e-39
	(b"00000000000111000010110010001010", b"00000000000000000000000000000000"),
	(b"10000000011000111010001110101111", b"10000000010001110111011100100101"), -- 2.58737e-39 + -9.15043e-39 = -6.56306e-39
	(b"00000000001000101101000111111111", b"00000000000000000000000000000000"),
	(b"00000000001101011100011011101011", b"00000000010110001001100011101010"), -- 3.19774e-39 + 4.93864e-39 = 8.13638e-39
	(b"00000000000101010001101001011111", b"00000000000000000000000000000000"),
	(b"00000000001001111000101110001011", b"00000000001111001010010111101010"), -- 1.93801e-39 + 3.63164e-39 = 5.56965e-39
	(b"10000000001000011010011111100110", b"00000000000000000000000000000000"),
	(b"00000000011100110011010101011100", b"00000000010100011000110101110110"), -- -3.0908e-39 + 1.05802e-38 = 7.48942e-39
	(b"00000000000011011110000001110000", b"00000000000000000000000000000000"),
	(b"10000000011111111001001001100111", b"10000000011100011011000111110111"), -- 1.27437e-39 + -1.17156e-38 = -1.04413e-38
	(b"00000000011001011000111001111100", b"00000000000000000000000000000000"),
	(b"10000000001011000011001111101010", b"00000000001110010101101010010010"), -- 9.3265e-39 + -4.05939e-39 = 5.26711e-39
	(b"00000000011101110011010100010000", b"00000000000000000000000000000000"),
	(b"00000000000110111000001011000110", b"00000000100100101011011111010110"), -- 1.09475e-38 + 2.52647e-39 = 1.34739e-38
	(b"00000000000011010001000001000100", b"00000000000000000000000000000000"),
	(b"00000000010011010101000011010101", b"00000000010110100110000100011001"), -- 1.1997e-39 + 7.10033e-39 = 8.30003e-39
	(b"00000000010011001010010110010010", b"00000000000000000000000000000000"),
	(b"10000000001100110101010101101100", b"00000000000110010101000000100110"), -- 7.03889e-39 + -4.71425e-39 = 2.32464e-39
	(b"10000000010111011010000000001111", b"00000000000000000000000000000000"),
	(b"10000000011101001100001111010011", b"10000000110100100110001111100010"), -- -8.59812e-39 + -1.07232e-38 = -1.93213e-38
	(b"00000000001100011001101010001111", b"00000000000000000000000000000000"),
	(b"10000000011101101010100000111101", b"10000000010001010000110110101110"), -- 4.55538e-39 + -1.08969e-38 = -6.34156e-39
	(b"10000000011110010111100110000101", b"00000000000000000000000000000000"),
	(b"10000000000001110101001000101111", b"10000000100000001100101110110100"), -- -1.11557e-38 + -6.7233e-40 = -1.1828e-38
	(b"00000000010000011100011101010010", b"00000000000000000000000000000000"),
	(b"00000000011101001100110001111000", b"00000000101101101001001111001010"), -- 6.04081e-39 + 1.07263e-38 = 1.67671e-38
	(b"10000000000101111111111011011001", b"00000000000000000000000000000000"),
	(b"10000000000101000000000001011001", b"10000000001010111111111100110010"), -- -2.20364e-39 + -1.83683e-39 = -4.04047e-39
	(b"10000000011100001000000001111000", b"00000000000000000000000000000000"),
	(b"10000000011110010111011100010110", b"10000000111010011111011110001110"), -- -1.03317e-38 + -1.11548e-38 = -2.14865e-38
	(b"00000000010110111010101110000011", b"00000000000000000000000000000000"),
	(b"10000000011000111101000011000000", b"10000000000010000010010100111101"), -- 8.41856e-39 + -9.1666e-39 = -7.48043e-40
	(b"10000000011000011100010110111011", b"00000000000000000000000000000000"),
	(b"00000000011100100001100100101000", b"00000000000100000101001101101101"), -- -8.97898e-39 + 1.04783e-38 = 1.4993e-39
	(b"00000000001110000001111001110010", b"00000000000000000000000000000000"),
	(b"00000000001000110101000111011111", b"00000000010110110111000001010001"), -- 5.15371e-39 + 3.24361e-39 = 8.39732e-39
	(b"10000000000100100111101111011000", b"00000000000000000000000000000000"),
	(b"00000000000000110101011101011100", b"10000000000011110010010001111100"), -- -1.69747e-39 + 3.06845e-40 = -1.39062e-39
	(b"00000000011010110000100010101000", b"00000000000000000000000000000000"),
	(b"10000000010100001000100110010011", b"00000000000110100111111100010101"), -- 9.8295e-39 + -7.39619e-39 = 2.43331e-39
	(b"00000000010011101111110001101000", b"00000000000000000000000000000000"),
	(b"00000000011010000111110100110010", b"00000000101101110111100110011010"), -- 7.25372e-39 + 9.5958e-39 = 1.68495e-38
	(b"00000000000011100100110110011110", b"00000000000000000000000000000000"),
	(b"00000000010011100110011000001100", b"00000000010111001011001110101010"), -- 1.31354e-39 + 7.19978e-39 = 8.51332e-39
	(b"10000000000110111010001010110110", b"00000000000000000000000000000000"),
	(b"10000000001001101100000001011111", b"10000000010000100110001100010101"), -- -2.53793e-39 + -3.55876e-39 = -6.09669e-39
	(b"10000000010000111110000011001000", b"00000000000000000000000000000000"),
	(b"10000000011001010000000101101001", b"10000000101010001110001000110001"), -- -6.23361e-39 + -9.27589e-39 = -1.55095e-38
	(b"10000000001000110000111111111110", b"00000000000000000000000000000000"),
	(b"00000000011010100011111100011100", b"00000000010001110010111100011110"), -- -3.21998e-39 + 9.7572e-39 = 6.53722e-39
	(b"00000000010001110110110111100011", b"00000000000000000000000000000000"),
	(b"00000000001111000110011000001010", b"00000000100000111101001111101101"), -- 6.55974e-39 + 5.54673e-39 = 1.21065e-38
	(b"00000000001001100100111010000010", b"00000000000000000000000000000000"),
	(b"10000000011010001111000100000110", b"10000000010000101010001010000100"), -- 3.51791e-39 + -9.63735e-39 = -6.11944e-39
	(b"00000000010011011110111011111001", b"00000000000000000000000000000000"),
	(b"00000000000001111010010101000001", b"00000000010101011001010000111010"), -- 7.15706e-39 + 7.0213e-40 = 7.85919e-39
	(b"10000000001110110011010010011110", b"00000000000000000000000000000000"),
	(b"10000000010100000110101111100111", b"10000000100010111010000010000101"), -- -5.43717e-39 + -7.38555e-39 = -1.28227e-38
	(b"00000000011101111010100010000000", b"00000000000000000000000000000000"),
	(b"10000000010000100101110000011100", b"00000000001101010100110001100100"), -- 1.09889e-38 + -6.09419e-39 = 4.89469e-39
	(b"00000000010111101001001110111011", b"00000000000000000000000000000000"),
	(b"00000000001111011000010100010110", b"00000000100111000001100011010001"), -- 8.68553e-39 + 5.64971e-39 = 1.43352e-38
	(b"10000000010101111010111110000100", b"00000000000000000000000000000000"),
	(b"10000000011001000111111110011110", b"10000000101111000010111100100010"), -- -8.05265e-39 + -9.22933e-39 = -1.7282e-38
	(b"10000000011000100111111101111001", b"00000000000000000000000000000000"),
	(b"10000000000001000110100100001101", b"10000000011001101110100010000110"), -- -9.04561e-39 + -4.05027e-40 = -9.45063e-39
	(b"00000000011000011100111001101000", b"00000000000000000000000000000000"),
	(b"00000000000010101010111101110110", b"00000000011011000111110111011110"), -- 8.98209e-39 + 9.81298e-40 = 9.96339e-39
	(b"00000000011011011110110101101011", b"00000000000000000000000000000000"),
	(b"00000000000111100011111111101101", b"00000000100011000010110101011000"), -- 1.00952e-38 + 2.778e-39 = 1.28732e-38
	(b"10000000000010110000011110110010", b"00000000000000000000000000000000"),
	(b"10000000010111111100001011111011", b"10000000011010101100101010101101"), -- -1.01295e-39 + -8.79432e-39 = -9.80727e-39
	(b"00000000011010000011010000111001", b"00000000000000000000000000000000"),
	(b"10000000011101011000001000110110", b"10000000000011010100110111111101"), -- 9.56963e-39 + -1.07915e-38 = -1.22184e-39
	(b"10000000010101010110111001011010", b"00000000000000000000000000000000"),
	(b"10000000011100010001010111011010", b"10000000110001101000010000110100"), -- -7.8456e-39 + -1.03852e-38 = -1.82309e-38
	(b"00000000000111010101100110101100", b"00000000000000000000000000000000"),
	(b"00000000011100110101010011100110", b"00000000100100001010111010010010"), -- 2.6954e-39 + 1.05915e-38 = 1.32869e-38
	(b"10000000001111011001001010000011", b"00000000000000000000000000000000"),
	(b"00000000011000100110100000111110", b"00000000001001001101010110111011"), -- -5.65452e-39 + 9.03727e-39 = 3.38275e-39
	(b"10000000011111111011011110000010", b"00000000000000000000000000000000"),
	(b"00000000010011111101101110011010", b"10000000001011111101101111101000"), -- -1.17289e-38 + 7.33378e-39 = -4.39516e-39
	(b"10000000001011001110010011001010", b"00000000000000000000000000000000"),
	(b"10000000011011111011101101000111", b"10000000100111001010000000010001"), -- -4.12284e-39 + -1.02609e-38 = -1.43838e-38
	(b"10000000010000000110101011111111", b"00000000000000000000000000000000"),
	(b"10000000011001011000001000011101", b"10000000101001011110110100011100"), -- -5.91585e-39 + -9.32206e-39 = -1.52379e-38
	(b"10000000001010000000111100111010", b"00000000000000000000000000000000"),
	(b"00000000011001010110011011100101", b"00000000001111010101011110101011"), -- -3.67888e-39 + 9.3123e-39 = 5.63341e-39
	(b"10000000011110010110011011101011", b"00000000000000000000000000000000"),
	(b"10000000000101001101001111111100", b"10000000100011100011101011100111"), -- -1.1149e-38 + -1.91276e-39 = -1.30618e-38
	(b"10000000001001000011111101010110", b"00000000000000000000000000000000"),
	(b"10000000001110101101100100010111", b"10000000010111110001100001101101"), -- -3.3288e-39 + -5.40434e-39 = -8.73313e-39
	(b"00000000001000011001011011100100", b"00000000000000000000000000000000"),
	(b"10000000010100110011011111111000", b"10000000001100011010000100010100"), -- 3.0847e-39 + -7.64242e-39 = -4.55772e-39
	(b"00000000001010000110110001001111", b"00000000000000000000000000000000"),
	(b"10000000001010110001111011011101", b"10000000000000101011001010001110"), -- 3.71227e-39 + -3.96e-39 = -2.47724e-40
	(b"10000000001111111011010101001010", b"00000000000000000000000000000000"),
	(b"00000000000110001100101111001000", b"10000000001001101110100110000010"), -- -5.85067e-39 + 2.27715e-39 = -3.57352e-39
	(b"00000000011100100010000100001111", b"00000000000000000000000000000000"),
	(b"10000000010000011100001010011000", b"00000000001100000101111001110111"), -- 1.04811e-38 + -6.03911e-39 = 4.44199e-39
	(b"00000000011100011100001011001011", b"00000000000000000000000000000000"),
	(b"10000000011001011001101001010000", b"00000000000011000010100001111011"), -- 1.04473e-38 + -9.33074e-39 = 1.11655e-39
	(b"10000000010100100000110101110000", b"00000000000000000000000000000000"),
	(b"10000000010100001101110001000101", b"10000000101000101110100110110101"), -- -7.53533e-39 + -7.42586e-39 = -1.49612e-38
	(b"10000000000000011101010111111010", b"00000000000000000000000000000000"),
	(b"10000000010101110001010100111010", b"10000000010110001110101100110100"), -- -1.68596e-40 + -7.9973e-39 = -8.1659e-39
	(b"00000000011011010100111101100010", b"00000000000000000000000000000000"),
	(b"00000000011110111000100010101000", b"00000000111010001101100000001010"), -- 1.00385e-38 + 1.13448e-38 = 2.13833e-38
	(b"00000000000010100101111101110101", b"00000000000000000000000000000000"),
	(b"00000000011101000001001000110011", b"00000000011111100111000110101000"), -- 9.52598e-40 + 1.06594e-38 = 1.1612e-38
	(b"10000000000001110100001100011100", b"00000000000000000000000000000000"),
	(b"00000000011010110010000110000010", b"00000000011000111101111001100110"), -- -6.66923e-40 + 9.83842e-39 = 9.1715e-39
	(b"10000000011000101010101011111010", b"00000000000000000000000000000000"),
	(b"10000000010110001000101011101101", b"10000000101110110011010111100111"), -- -9.06121e-39 + -8.13136e-39 = -1.71926e-38
	(b"10000000000001101111101000100111", b"00000000000000000000000000000000"),
	(b"10000000001101111011010010001111", b"10000000001111101010111010110110"), -- -6.40751e-40 + -5.11572e-39 = -5.75648e-39
	(b"10000000000101000110101010010100", b"00000000000000000000000000000000"),
	(b"00000000001110100110110100011001", b"00000000001001100000001010000101"), -- -1.87494e-39 + 5.3656e-39 = 3.49065e-39
	(b"00000000010000001001001111101111", b"00000000000000000000000000000000"),
	(b"10000000000001111110111011011000", b"00000000001110001010010100010111"), -- 5.93054e-39 + -7.28529e-40 = 5.20201e-39
	(b"00000000010010101111001100110001", b"00000000000000000000000000000000"),
	(b"10000000001100100001111010011010", b"00000000000110001101010010010111"), -- 6.88307e-39 + -4.60275e-39 = 2.28031e-39
	(b"10000000001011011101000110100111", b"00000000000000000000000000000000"),
	(b"00000000001101010011001101101001", b"00000000000001110110000111000010"), -- -4.20781e-39 + 4.88572e-39 = 6.77917e-40
	(b"10000000001011010011101111000011", b"00000000000000000000000000000000"),
	(b"10000000000111000101001101001011", b"10000000010010011000111100001110"), -- -4.15404e-39 + -2.60127e-39 = -6.75531e-39
	(b"00000000010110010000000101111100", b"00000000000000000000000000000000"),
	(b"00000000010111001110101010110101", b"00000000101101011110110000110001"), -- 8.17389e-39 + 8.53306e-39 = 1.6707e-38
	(b"10000000001100000111101010111100", b"00000000000000000000000000000000"),
	(b"10000000011101100111000010100110", b"10000000101001101110101101100010"), -- -4.45213e-39 + -1.0877e-38 = -1.53291e-38
	(b"00000000010010010110110100111011", b"00000000000000000000000000000000"),
	(b"10000000001010101111101101011001", b"00000000000111100111000111100010"), -- 6.74318e-39 + -3.94726e-39 = 2.79592e-39
	(b"10000000000110111001100010010110", b"00000000000000000000000000000000"),
	(b"00000000001001110001011100000110", b"00000000000010110111111001110000"), -- -2.5343e-39 + 3.58984e-39 = 1.05555e-39
	(b"10000000001111100110111111010010", b"00000000000000000000000000000000"),
	(b"10000000001100000000011110001010", b"10000000011011100111011101011100"), -- -5.73391e-39 + -4.41081e-39 = -1.01447e-38
	(b"10000000010001010001110011101000", b"00000000000000000000000000000000"),
	(b"10000000010011000000101011101101", b"10000000100100010010011111010101"), -- -6.34702e-39 + -6.98342e-39 = -1.33304e-38
	(b"00000000011011010110100011010010", b"00000000000000000000000000000000"),
	(b"00000000001101100100010001010101", b"00000000101000111010110100100111"), -- 1.00477e-38 + 4.98363e-39 = 1.50313e-38
	(b"10000000000100000100000011010001", b"00000000000000000000000000000000"),
	(b"00000000001001110000011000011011", b"00000000000101101100010101001010"), -- -1.49262e-39 + 3.58377e-39 = 2.09115e-39
	(b"00000000010111110011010100110010", b"00000000000000000000000000000000"),
	(b"00000000011010101000000110001111", b"00000000110010011011011011000001"), -- 8.74346e-39 + 9.78104e-39 = 1.85245e-38
	(b"10000000000001011000100111010110", b"00000000000000000000000000000000"),
	(b"00000000001000010100111001001101", b"00000000000110111100010001110111"), -- -5.08624e-40 + 3.05866e-39 = 2.55004e-39
	(b"00000000011011011000111011101110", b"00000000000000000000000000000000"),
	(b"00000000011110101010101001100110", b"00000000111010000011100101010100"), -- 1.00613e-38 + 1.12651e-38 = 2.13264e-38
	(b"10000000000101111001111011110011", b"00000000000000000000000000000000"),
	(b"00000000000100111011000011100110", b"10000000000000111110111000001101"), -- -2.16924e-39 + 1.80833e-39 = -3.60903e-40
	(b"00000000000110000110100110000110", b"00000000000000000000000000000000"),
	(b"00000000011111101001100111101011", b"00000000100101110000001101110001"), -- 2.24191e-39 + 1.16265e-38 = 1.38684e-38
	(b"10000000000101100001111001110000", b"00000000000000000000000000000000"),
	(b"10000000001000100111111111000010", b"10000000001110001001111000110010"), -- -2.0313e-39 + -3.16824e-39 = -5.19954e-39
	(b"00000000011001110011010111100111", b"00000000000000000000000000000000"),
	(b"10000000010101001010101000001101", b"00000000000100101000101111011010"), -- 9.47839e-39 + -7.77518e-39 = 1.70321e-39
	(b"10000000000011001011000101110010", b"00000000000000000000000000000000"),
	(b"00000000001111001101111100111110", b"00000000001100000010110111001100"), -- -1.16568e-39 + 5.59021e-39 = 4.42453e-39
	(b"00000000010100000001101111000100", b"00000000000000000000000000000000"),
	(b"00000000010010111111111110000111", b"00000000100111000001101101001011"), -- 7.3568e-39 + 6.97933e-39 = 1.43361e-38
	(b"10000000000010001111111110010110", b"00000000000000000000000000000000"),
	(b"00000000011111000111110101010110", b"00000000011100110111110111000000"), -- -8.26371e-40 + 1.14326e-38 = 1.06062e-38
	(b"00000000001011000100100100011011", b"00000000000000000000000000000000"),
	(b"00000000001101011011011001111110", b"00000000011000011111111110011001"), -- 4.06699e-39 + 4.93275e-39 = 8.99973e-39
	(b"10000000010000001110100111101000", b"00000000000000000000000000000000"),
	(b"10000000010010010001111011001000", b"10000000100010100000100010110000"), -- -5.96138e-39 + -6.71503e-39 = -1.26764e-38
	(b"10000000000010101101101011110100", b"00000000000000000000000000000000"),
	(b"10000000000010000101101001100100", b"10000000000100110011010101011000"), -- -9.96901e-40 + -7.6711e-40 = -1.76401e-39
	(b"00000000000101000011111001010001", b"00000000000000000000000000000000"),
	(b"10000000010010001110001111000100", b"10000000001101001010010101110011"), -- 1.85906e-39 + -6.69386e-39 = -4.8348e-39
	(b"10000000011011100011101011001010", b"00000000000000000000000000000000"),
	(b"10000000001001100011100111101100", b"10000000100101000111010010110110"), -- -1.0123e-38 + -3.51053e-39 = -1.36335e-38
	(b"10000000011001001110101010000100", b"00000000000000000000000000000000"),
	(b"10000000001011000010000110111100", b"10000000100100010000110001000000"), -- -9.26768e-39 + -4.05286e-39 = -1.33205e-38
	(b"00000000000011010000010100001011", b"00000000000000000000000000000000"),
	(b"10000000000100000111110111111100", b"10000000000000110111100011110001"), -- 1.19567e-39 + -1.51456e-39 = -3.18892e-40
	(b"10000000001000001010110111001101", b"00000000000000000000000000000000"),
	(b"10000000000010011001111101101011", b"10000000001010100100110100111000"), -- -3.00108e-39 + -8.83708e-40 = -3.88479e-39
	(b"10000000000110000101110100011111", b"00000000000000000000000000000000"),
	(b"10000000001000101001001111110011", b"10000000001110101111000100010010"), -- -2.23746e-39 + -3.17548e-39 = -5.41294e-39
	(b"00000000011110011100111101110000", b"00000000000000000000000000000000"),
	(b"10000000011001101010111000011011", b"00000000000100110010000101010101"), -- 1.11865e-38 + -9.42968e-39 = 1.75683e-39
	(b"00000000000001110001001000000010", b"00000000000000000000000000000000"),
	(b"10000000000100100011111101101111", b"10000000000010110010110101101101"), -- 6.49308e-40 + -1.67579e-39 = -1.02649e-39
	(b"00000000010010011000110000011100", b"00000000000000000000000000000000"),
	(b"00000000010111010011001010111011", b"00000000101001101011111011010111"), -- 6.75425e-39 + 8.5589e-39 = 1.53132e-38
	(b"10000000010111010010110111110101", b"00000000000000000000000000000000"),
	(b"10000000001001010011011110111111", b"10000000100000100110010110110100"), -- -8.55719e-39 + -3.41791e-39 = -1.19751e-38
	(b"00000000011100101001011010011000", b"00000000000000000000000000000000"),
	(b"10000000011100011011010111101101", b"00000000000000001110000010101011"), -- 1.05233e-38 + -1.04427e-38 = 8.05957e-41
	(b"10000000011000011100011110001101", b"00000000000000000000000000000000"),
	(b"00000000001001010111001111101110", b"10000000001111000101001110011111"), -- -8.97963e-39 + 3.4395e-39 = -5.54013e-39
	(b"00000000011010000111100100110111", b"00000000000000000000000000000000"),
	(b"00000000010100000101001100101001", b"00000000101110001100110001100000"), -- 9.59438e-39 + 7.37667e-39 = 1.6971e-38
	(b"00000000010011101101101010011011", b"00000000000000000000000000000000"),
	(b"00000000011101010111001101000010", b"00000000110001000100110111011101"), -- 7.24159e-39 + 1.07861e-38 = 1.80277e-38
	(b"00000000000001010111011000101001", b"00000000000000000000000000000000"),
	(b"00000000000101100011110101000100", b"00000000000110111011001101101101"), -- 5.01565e-40 + 2.04236e-39 = 2.54392e-39
	(b"10000000001100100110110010011100", b"00000000000000000000000000000000"),
	(b"10000000000010101010001000001111", b"10000000001111010000111010101011"), -- -4.63074e-39 + -9.76491e-40 = -5.60723e-39
	(b"10000000000110000011100010101101", b"00000000000000000000000000000000"),
	(b"10000000010110001010010010101101", b"10000000011100001101110101011010"), -- -2.22438e-39 + -8.1406e-39 = -1.0365e-38
	(b"10000000000101110000011010100100", b"00000000000000000000000000000000"),
	(b"00000000011100111001011111000011", b"00000000010111001001000100011111"), -- -2.1146e-39 + 1.06155e-38 = 8.50093e-39
	(b"00000000000011000010110110001111", b"00000000000000000000000000000000"),
	(b"00000000011111101000110000100000", b"00000000100010101011100110101111"), -- 1.11837e-39 + 1.16215e-38 = 1.27399e-38
	(b"00000000000110110101111110011111", b"00000000000000000000000000000000"),
	(b"10000000011111000011001000011000", b"10000000011000001101001001111001"), -- 2.51386e-39 + -1.14056e-38 = -8.89171e-39
	(b"00000000010001000101011010110101", b"00000000000000000000000000000000"),
	(b"10000000001000001001010000100110", b"00000000001000111100001010001111"), -- 6.27592e-39 + -2.99188e-39 = 3.28404e-39
	(b"10000000001110111110111100001111", b"00000000000000000000000000000000"),
	(b"00000000011000001010100001101100", b"00000000001001001011100101011101"), -- -5.50405e-39 + 8.87663e-39 = 3.37257e-39
	(b"00000000010111100101010111000100", b"00000000000000000000000000000000"),
	(b"10000000001000000110101101000011", b"00000000001111011110101010000001"), -- 8.6633e-39 + -2.97721e-39 = 5.68609e-39
	(b"10000000000000011000110100011110", b"00000000000000000000000000000000"),
	(b"10000000001000010001000110010001", b"10000000001000101001111010101111"), -- -1.42459e-40 + -3.03687e-39 = -3.17933e-39
	(b"10000000000000010010100001001110", b"00000000000000000000000000000000"),
	(b"00000000010101011010000110000101", b"00000000010101000111100100110111"), -- -1.06294e-40 + 7.86396e-39 = 7.75767e-39
	(b"10000000000001110010111101111011", b"00000000000000000000000000000000"),
	(b"10000000010010010101111111101111", b"10000000010100001000111101101010"), -- -6.59881e-40 + -6.73841e-39 = -7.39829e-39
	(b"10000000011100110011000011010111", b"00000000000000000000000000000000"),
	(b"10000000000101111100010110000011", b"10000000100010101111011001011010"), -- -1.05786e-38 + -2.18307e-39 = -1.27617e-38
	(b"00000000010110101100101100001111", b"00000000000000000000000000000000"),
	(b"00000000011001100111001010101001", b"00000000110000010011110110111000"), -- 8.33804e-39 + 9.40835e-39 = 1.77464e-38
	(b"10000000010101111101000111011100", b"00000000000000000000000000000000"),
	(b"00000000001101110010011011111101", b"10000000001000001010101011011111"), -- -8.06497e-39 + 5.06494e-39 = -3.00003e-39
	(b"00000000000001111100010011010011", b"00000000000000000000000000000000"),
	(b"10000000000001010100000101010011", b"00000000000000101000001110000000"), -- 7.13456e-40 + -4.82611e-40 = 2.30844e-40
	(b"00000000000001100010000101001011", b"00000000000000000000000000000000"),
	(b"10000000001110110100001110110100", b"10000000001101010010001001101001"), -- 5.62956e-40 + -5.44258e-39 = -4.87963e-39
	(b"00000000010011111111011001011111", b"00000000000000000000000000000000"),
	(b"10000000000101011111001000001011", b"00000000001110100000010001010100"), -- 7.34339e-39 + -2.01537e-39 = 5.32801e-39
	(b"10000000010111101110101000010110", b"00000000000000000000000000000000"),
	(b"10000000000110000010110100000011", b"10000000011101110001011100011001"), -- -8.71651e-39 + -2.2202e-39 = -1.09367e-38
	(b"00000000010010111111011000010001", b"00000000000000000000000000000000"),
	(b"00000000000000100101101101111011", b"00000000010011100101000110001100"), -- 6.97593e-39 + 2.16488e-40 = 7.19242e-39
	(b"10000000000000100000011101101000", b"00000000000000000000000000000000"),
	(b"00000000010110011010001010110100", b"00000000010101111001101101001100"), -- -1.86328e-40 + 8.23173e-39 = 8.0454e-39
	(b"00000000000111011110101010100011", b"00000000000000000000000000000000"),
	(b"10000000011010010001111010000100", b"10000000010010110011001111100001"), -- 2.7474e-39 + -9.65367e-39 = -6.90627e-39
	(b"10000000000010100011011110011010", b"00000000000000000000000000000000"),
	(b"10000000011101011110101101000101", b"10000000100000000010001011011111"), -- -9.38301e-40 + -1.08292e-38 = -1.17675e-38
	(b"00000000011000101111011011010011", b"00000000000000000000000000000000"),
	(b"10000000000011101111101011101001", b"00000000010100111111101111101010"), -- 9.08842e-39 + -1.37571e-39 = 7.71272e-39
	(b"10000000010010000101001001010110", b"00000000000000000000000000000000"),
	(b"00000000000011111100110101001111", b"10000000001110001000010100000111"), -- -6.64169e-39 + 1.45118e-39 = -5.19051e-39
	(b"00000000000010111111000000001001", b"00000000000000000000000000000000"),
	(b"00000000001000010011110001100100", b"00000000001011010010110001101101"), -- 1.0963e-39 + 3.05224e-39 = 4.14853e-39
	(b"10000000001010001111111000111010", b"00000000000000000000000000000000"),
	(b"10000000000111010101100011011011", b"10000000010001100101011100010101"), -- -3.76462e-39 + -2.6951e-39 = -6.45972e-39
	(b"10000000000101100011011110011000", b"00000000000000000000000000000000"),
	(b"10000000000010110110110011011100", b"10000000001000011010010001110100"), -- -2.04032e-39 + -1.04924e-39 = -3.08957e-39
	(b"00000000010101100001101011100001", b"00000000000000000000000000000000"),
	(b"10000000011110011111101110001100", b"10000000001000111110000010101011"), -- 7.9075e-39 + -1.12023e-38 = -3.29484e-39
	(b"10000000000001111111010110000010", b"00000000000000000000000000000000"),
	(b"10000000010001010110111101000000", b"10000000010011010110010011000010"), -- -7.3092e-40 + -6.37656e-39 = -7.10748e-39
	(b"00000000001000111000100011110111", b"00000000000000000000000000000000"),
	(b"00000000010100000110110101011010", b"00000000011100111111011001010001"), -- 3.26338e-39 + 7.38607e-39 = 1.06494e-38
	(b"00000000000001111000011100111100", b"00000000000000000000000000000000"),
	(b"10000000000000101010101101001110", b"00000000000001001101101111101110"), -- 6.91361e-40 + -2.45124e-40 = 4.46238e-40
	(b"00000000010111010000001000001001", b"00000000000000000000000000000000"),
	(b"00000000010111010001101110101001", b"00000000101110100001110110110010"), -- 8.54143e-39 + 8.55062e-39 = 1.70921e-38
	(b"10000000011010100001010001110100", b"00000000000000000000000000000000"),
	(b"00000000001000111001111101110000", b"10000000010001100111010100000100"), -- -9.7419e-39 + 3.27144e-39 = -6.47046e-39
	(b"00000000001000111010010011101110", b"00000000000000000000000000000000"),
	(b"10000000001110101111110011000011", b"10000000000101110101011111010101"), -- 3.27341e-39 + -5.41713e-39 = -2.14372e-39
	(b"00000000001000010000111100001000", b"00000000000000000000000000000000"),
	(b"00000000010011110011000100101111", b"00000000011100000100000000110111"), -- 3.03596e-39 + 7.27265e-39 = 1.03086e-38
	(b"10000000001001101000011100111110", b"00000000000000000000000000000000"),
	(b"00000000000100111101010001000111", b"10000000000100101011001011110111"), -- -3.53826e-39 + 1.82103e-39 = -1.71724e-39
	(b"10000000011000111100111100001011", b"00000000000000000000000000000000"),
	(b"00000000011010010111011100101100", b"00000000000001011010100000100001"), -- -9.16599e-39 + 9.68548e-39 = 5.19491e-40
	(b"00000000010101111111100000100001", b"00000000000000000000000000000000"),
	(b"00000000001100101101000110111110", b"00000000100010101100100111011111"), -- 8.0787e-39 + 4.66702e-39 = 1.27457e-38
	(b"10000000000110000101010110010101", b"00000000000000000000000000000000"),
	(b"10000000000011010011100101011101", b"10000000001001011000111011110010"), -- -2.23475e-39 + -1.21444e-39 = -3.44919e-39
	(b"10000000010110000111101100100111", b"00000000000000000000000000000000"),
	(b"00000000011100010101111101110001", b"00000000000110001110010001001010"), -- -8.1257e-39 + 1.04116e-38 = 2.28595e-39
	(b"00000000000011111111000101101100", b"00000000000000000000000000000000"),
	(b"00000000011110001110001010110101", b"00000000100010001101010000100001"), -- 1.46414e-39 + 1.11016e-38 = 1.25657e-38
	(b"00000000001000110000100110010101", b"00000000000000000000000000000000"),
	(b"00000000000110110101110100101001", b"00000000001111100110011010111110"), -- 3.21768e-39 + 2.51298e-39 = 5.73066e-39
	(b"00000000010010000110001110110011", b"00000000000000000000000000000000"),
	(b"10000000010001101011110001101001", b"00000000000000011010011101001010"), -- 6.64792e-39 + -6.49607e-39 = 1.51848e-40
	(b"10000000010110001000000101001010", b"00000000000000000000000000000000"),
	(b"00000000000011111111111000010100", b"10000000010010001000001100110110"), -- -8.1279e-39 + 1.46868e-39 = -6.65923e-39
	(b"10000000010100010011101011010001", b"00000000000000000000000000000000"),
	(b"10000000001011111010011111100011", b"10000000100000001110001010110100"), -- -7.45977e-39 + -4.37649e-39 = -1.18363e-38
	(b"00000000010001010111101110011001", b"00000000000000000000000000000000"),
	(b"10000000001001110101001001110010", b"00000000000111100010100100100111"), -- 6.38099e-39 + -3.61116e-39 = 2.76983e-39
	(b"10000000010100100110111100011010", b"00000000000000000000000000000000"),
	(b"00000000001011011111110010011110", b"10000000001001000111001001111100"), -- -7.57037e-39 + 4.22322e-39 = -3.34715e-39
	(b"10000000010010100011110010111001", b"00000000000000000000000000000000"),
	(b"10000000000001111101101011111110", b"10000000010100100001011110110111"), -- -6.81761e-39 + -7.21408e-40 = -7.53902e-39
	(b"10000000011111011110001100100011", b"00000000000000000000000000000000"),
	(b"10000000001000001100100010001101", b"10000000100111101010101110110000"), -- -1.15609e-38 + -3.01068e-39 = -1.45716e-38
	(b"00000000011011100001111000110111", b"00000000000000000000000000000000"),
	(b"00000000011111010000101000011001", b"00000000111010110010100001010000"), -- 1.01127e-38 + 1.14831e-38 = 2.15958e-38
	(b"00000000011001110101100001010111", b"00000000000000000000000000000000"),
	(b"00000000011101100111110110111110", b"00000000110111011101011000010101"), -- 9.49075e-39 + 1.08817e-38 = 2.03724e-38
	(b"00000000010000011100110000000110", b"00000000000000000000000000000000"),
	(b"10000000000000001011110111100011", b"00000000010000010000111000100011"), -- 6.0425e-39 + -6.81185e-41 = 5.97438e-39
	(b"00000000000011011101010011110110", b"00000000000000000000000000000000"),
	(b"10000000010111000111001101100001", b"10000000010011101001111001101011"), -- 1.27026e-39 + -8.49026e-39 = -7.22e-39
	(b"00000000010111010011000001000101", b"00000000000000000000000000000000"),
	(b"00000000010001001111001001011000", b"00000000101000100010001010011101"), -- 8.55802e-39 + 6.33175e-39 = 1.48898e-38
	(b"00000000000101000110111100010110", b"00000000000000000000000000000000"),
	(b"00000000011000111100110000001110", b"00000000011110000011101100100100"), -- 1.87656e-39 + 9.16492e-39 = 1.10415e-38
	(b"10000000011010111010011011100001", b"00000000000000000000000000000000"),
	(b"10000000010010100100110111110101", b"10000000101101011111010011010110"), -- -9.88626e-39 + -6.82379e-39 = -1.67101e-38
	(b"00000000010101000100001011000110", b"00000000000000000000000000000000"),
	(b"10000000000100110100101010000100", b"00000000010000001111100001000010"), -- 7.73814e-39 + -1.77161e-39 = 5.96653e-39
	(b"10000000011001000101000001101101", b"00000000000000000000000000000000"),
	(b"10000000000001101110011011010110", b"10000000011010110011011101000011"), -- -9.2124e-39 + -6.33821e-40 = -9.84622e-39
	(b"00000000001110111011110000111010", b"00000000000000000000000000000000"),
	(b"10000000010000000001001001110101", b"10000000000001000101011000111011"), -- 5.48582e-39 + -5.88409e-39 = -3.98276e-40
	(b"00000000000000101100000111000011", b"00000000000000000000000000000000"),
	(b"10000000011110101100000101000100", b"10000000011101111111111110000001"), -- 2.5318e-40 + -1.12733e-38 = -1.10201e-38
	(b"10000000001011111011000101011110", b"00000000000000000000000000000000"),
	(b"00000000000010001010000000001100", b"10000000001001110001000101010010"), -- -4.3799e-39 + 7.92098e-40 = -3.5878e-39
	(b"00000000000101110101110110110010", b"00000000000000000000000000000000"),
	(b"00000000011100011010111100100000", b"00000000100010010000110011010010"), -- 2.14583e-39 + 1.04402e-38 = 1.25861e-38
	(b"00000000011110000001000011000111", b"00000000000000000000000000000000"),
	(b"00000000001101000100101010110110", b"00000000101011000101101101111101"), -- 1.10263e-38 + 4.80225e-39 = 1.58285e-38
	(b"00000000000101001010011011010000", b"00000000000000000000000000000000"),
	(b"10000000011000001101001001100011", b"10000000010011000010101110010011"), -- 1.89655e-39 + -8.89168e-39 = -6.99513e-39
	(b"00000000010101110101010010000101", b"00000000000000000000000000000000"),
	(b"10000000010111110000111010101001", b"10000000000001111011101000100100"), -- 8.02001e-39 + -8.72963e-39 = -7.09623e-40
	(b"10000000001000011001100010101011", b"00000000000000000000000000000000"),
	(b"00000000000100101010001100011010", b"10000000000011101111010110010001"), -- -3.08534e-39 + 1.71155e-39 = -1.37379e-39
	(b"10000000001100111111100111001010", b"00000000000000000000000000000000"),
	(b"00000000001111101110000001110100", b"00000000000010101110011010101010"), -- -4.77322e-39 + 5.77432e-39 = 1.0011e-39
	(b"10000000000001101111100000100000", b"00000000000000000000000000000000"),
	(b"10000000001101110010101111111111", b"10000000001111100010010000011111"), -- -6.40023e-40 + -5.06674e-39 = -5.70676e-39
	(b"10000000010110010010001010000011", b"00000000000000000000000000000000"),
	(b"10000000011111000001011000010110", b"10000000110101010011100010011001"), -- -8.18574e-39 + -1.13955e-38 = -1.95813e-38
	(b"10000000010101111100101100101110", b"00000000000000000000000000000000"),
	(b"10000000001000011011101100011001", b"10000000011110011000011001000111"), -- -8.06258e-39 + -3.09769e-39 = -1.11603e-38
	(b"00000000001001110101010111010011", b"00000000000000000000000000000000"),
	(b"00000000001110110001010101100010", b"00000000011000100110101100110101"), -- 3.61237e-39 + 5.42596e-39 = 9.03834e-39
	(b"10000000000000011110111100011110", b"00000000000000000000000000000000"),
	(b"10000000010011101100000111101001", b"10000000010100001011000100000111"), -- -1.77615e-40 + -7.23273e-39 = -7.41035e-39
	(b"00000000010001100100111001000111", b"00000000000000000000000000000000"),
	(b"10000000011001111010100101011000", b"10000000001000010101101100010001"), -- 6.45657e-39 + -9.51981e-39 = -3.06324e-39
	(b"00000000001001011011001010010010", b"00000000000000000000000000000000"),
	(b"00000000001010011111101011110000", b"00000000010011111010110110000010"), -- 3.46197e-39 + 3.85527e-39 = 7.31725e-39
	(b"10000000000001101110010111011111", b"00000000000000000000000000000000"),
	(b"10000000001111001101010100001011", b"10000000010000111011101011101010"), -- -6.33475e-40 + -5.58656e-39 = -6.22003e-39
	(b"00000000000111100000101111001100", b"00000000000000000000000000000000"),
	(b"10000000001011100011000010101000", b"10000000000100000010010011011100"), -- 2.7593e-39 + -4.24189e-39 = -1.48259e-39
	(b"00000000001101010101000111111101", b"00000000000000000000000000000000"),
	(b"00000000011100000011100100001001", b"00000000101001011000101100000110"), -- 4.89669e-39 + 1.0306e-38 = 1.52027e-38
	(b"00000000011110110111110111010101", b"00000000000000000000000000000000"),
	(b"00000000011111011010111010011110", b"00000000111110010010110001110011"), -- 1.13409e-38 + 1.15421e-38 = 2.2883e-38
	(b"00000000011110101001111000010110", b"00000000000000000000000000000000"),
	(b"00000000010001110010101110010011", b"00000000110000011100100110101001"), -- 1.12606e-38 + 6.53595e-39 = 1.77966e-38
	(b"10000000001101101101001010111101", b"00000000000000000000000000000000"),
	(b"10000000011011000000111101111111", b"10000000101000101110001000111100"), -- -5.03472e-39 + -9.92379e-39 = -1.49585e-38
	(b"00000000010001001000100010011101", b"00000000000000000000000000000000"),
	(b"00000000001110101110110101100010", b"00000000011111110111010111111111"), -- 6.29382e-39 + 5.41162e-39 = 1.17054e-38
	(b"10000000011011111000100100001010", b"00000000000000000000000000000000"),
	(b"00000000001000010101111001000010", b"10000000010011100010101011001000"), -- -1.02429e-38 + 3.06438e-39 = -7.17852e-39
	(b"00000000001110000010010100110010", b"00000000000000000000000000000000"),
	(b"00000000001111011011110011010110", b"00000000011101011110001000001000"), -- 5.15613e-39 + 5.66971e-39 = 1.08258e-38
	(b"00000000011111011110110111011011", b"00000000000000000000000000000000"),
	(b"00000000011100110100011110011011", b"00000000111100010011010101110110"), -- 1.15648e-38 + 1.05868e-38 = 2.21515e-38
	(b"10000000001100010010110000011111", b"00000000000000000000000000000000"),
	(b"00000000011100011100101000100010", b"00000000010000001001111000000011"), -- -4.51577e-39 + 1.04499e-38 = 5.93416e-39
	(b"10000000011010011010110010101000", b"00000000000000000000000000000000"),
	(b"10000000010101000110101001101001", b"10000000101111100001011100010001"), -- -9.70466e-39 + -7.75235e-39 = -1.7457e-38
	(b"00000000011011111101111111011010", b"00000000000000000000000000000000"),
	(b"00000000001111100011111101100000", b"00000000101011100001111100111010"), -- 1.0274e-38 + 5.71654e-39 = 1.59906e-38
	(b"10000000001110110000110000111101", b"00000000000000000000000000000000"),
	(b"10000000011111001000000000100100", b"10000000101101111000110001100001"), -- -5.42268e-39 + -1.14336e-38 = -1.68563e-38
	(b"10000000011100110000000101101001", b"00000000000000000000000000000000"),
	(b"00000000010000000101000111100000", b"10000000001100101010111110001001"), -- -1.05616e-38 + 5.90684e-39 = -4.65474e-39
	(b"10000000001100101001100011000111", b"00000000000000000000000000000000"),
	(b"10000000011011010010110010001100", b"10000000100111111100010101010011"), -- -4.64658e-39 + -1.0026e-38 = -1.46726e-38
	(b"00000000010101000010100110110110", b"00000000000000000000000000000000"),
	(b"00000000010110000000101010100110", b"00000000101011000011010001011100"), -- 7.72914e-39 + 8.08534e-39 = 1.58145e-38
	(b"10000000000011011001010011011000", b"00000000000000000000000000000000"),
	(b"10000000001001010000001010100100", b"10000000001100101001011101111100"), -- -1.24726e-39 + -3.39886e-39 = -4.64612e-39
	(b"00000000010010001101100111100110", b"00000000000000000000000000000000"),
	(b"10000000001110111111101101101000", b"00000000000011001101111001111110"), -- 6.69032e-39 + -5.50848e-39 = 1.18184e-39
	(b"10000000010110000101010100101001", b"00000000000000000000000000000000"),
	(b"10000000010111000101110100111111", b"10000000101101001011001001101000"), -- -8.11207e-39 + -8.48232e-39 = -1.65944e-38
	(b"10000000000010111010101101011100", b"00000000000000000000000000000000"),
	(b"10000000010110010011001000101110", b"10000000011001001101110110001010"), -- -1.07166e-39 + -8.19136e-39 = -9.26302e-39
	(b"00000000001001000010110100111000", b"00000000000000000000000000000000"),
	(b"10000000011011011100011101101001", b"10000000010010011001101000110001"), -- 3.3223e-39 + -1.00816e-38 = -6.7593e-39
	(b"10000000011001011100101000100000", b"00000000000000000000000000000000"),
	(b"00000000011011100000110111101001", b"00000000000010000100001111001001"), -- -9.34789e-39 + 1.01069e-38 = 7.59001e-40
	(b"10000000010110011100001011011100", b"00000000000000000000000000000000"),
	(b"00000000010110101111011011011111", b"00000000000000010011010000000011"), -- -8.24326e-39 + 8.35376e-39 = 1.10494e-40
	(b"00000000011100001000111000010001", b"00000000000000000000000000000000"),
	(b"10000000000111000101100001101100", b"00000000010101000011010110100101"), -- 1.03365e-38 + -2.60311e-39 = 7.73343e-39
	(b"00000000001000100111111111011011", b"00000000000000000000000000000000"),
	(b"10000000000011011100111111100110", b"00000000000101001010111111110101"), -- 3.16827e-39 + -1.26844e-39 = 1.89983e-39
	(b"10000000011010011010010011110101", b"00000000000000000000000000000000"),
	(b"00000000011010010001011011110101", b"10000000000000001000111000000000"), -- -9.7019e-39 + 9.65096e-39 = -5.094e-41
	(b"10000000001110011000000100100000", b"00000000000000000000000000000000"),
	(b"00000000010110100100111101101010", b"00000000001000001100111001001010"), -- -5.28094e-39 + 8.29368e-39 = 3.01274e-39
	(b"10000000000101111011100010100110", b"00000000000000000000000000000000"),
	(b"10000000001111101010100101011111", b"10000000010101100110001000000101"), -- -2.17846e-39 + -5.75456e-39 = -7.93302e-39
	(b"10000000001011100100011010100001", b"00000000000000000000000000000000"),
	(b"10000000001001100011101101111010", b"10000000010101001000001000011011"), -- -4.24977e-39 + -3.51109e-39 = -7.76085e-39
	(b"00000000011111101111000011100010", b"00000000000000000000000000000000"),
	(b"10000000010010101101000101110110", b"00000000001101000001111101101100"), -- 1.16577e-38 + -6.87097e-39 = 4.78672e-39
	(b"10000000000100011110010110101011", b"00000000000000000000000000000000"),
	(b"10000000001010100111101111100000", b"10000000001111000110000110001011"), -- -1.64359e-39 + -3.90153e-39 = -5.54512e-39
	(b"10000000010110001100001011110110", b"00000000000000000000000000000000"),
	(b"10000000000101110100111100100001", b"10000000011100000001001000010111"), -- -8.15146e-39 + -2.1406e-39 = -1.02921e-38
	(b"00000000010000100001000000011110", b"00000000000000000000000000000000"),
	(b"10000000001101100101000111011110", b"00000000000010111011111001000000"), -- 6.06692e-39 + -4.98849e-39 = 1.07844e-39
	(b"10000000001010100100110101110001", b"00000000000000000000000000000000"),
	(b"10000000010001010001001001010111", b"10000000011011110101111111001000"), -- -3.88487e-39 + -6.34323e-39 = -1.02281e-38
	(b"10000000001011000110100101100010", b"00000000000000000000000000000000"),
	(b"00000000000010000000110111011100", b"10000000001001000101101110000110"), -- -4.07857e-39 + 7.39656e-40 = -3.33891e-39
	(b"10000000000001110000111001101111", b"00000000000000000000000000000000"),
	(b"10000000011111101101001010010011", b"10000000100001011110000100000010"), -- -6.48026e-40 + -1.16468e-38 = -1.22948e-38
	(b"00000000010000000100110110101110", b"00000000000000000000000000000000"),
	(b"00000000010010100010111001001101", b"00000000100010100111101111111011"), -- 5.90534e-39 + 6.81244e-39 = 1.27178e-38
	(b"10000000010001100001000011011010", b"00000000000000000000000000000000"),
	(b"00000000011100001111110111100011", b"00000000001010101110110100001001"), -- -6.43453e-39 + 1.03767e-38 = 3.94212e-39
	(b"00000000001001110000101001111010", b"00000000000000000000000000000000"),
	(b"10000000011111110110011110111001", b"10000000010110000101110100111111"), -- 3.58534e-39 + -1.17003e-38 = -8.11497e-39
	(b"00000000011110101011111101100000", b"00000000000000000000000000000000"),
	(b"10000000000000010011010010111111", b"00000000011110011000101010100001"), -- 1.12726e-38 + -1.10757e-40 = 1.11618e-38
	(b"00000000011100000001011100101011", b"00000000000000000000000000000000"),
	(b"00000000000010100111100010001111", b"00000000011110101000111110111010"), -- 1.02939e-38 + 9.61603e-40 = 1.12555e-38
	(b"00000000000011010101110111110100", b"00000000000000000000000000000000"),
	(b"00000000011101011110001111100101", b"00000000100000110100000111011001"), -- 1.22757e-39 + 1.08265e-38 = 1.20541e-38
	(b"10000000001100111001110010010110", b"00000000000000000000000000000000"),
	(b"10000000011001110011001111010001", b"10000000100110101101000001100111"), -- -4.73978e-39 + -9.47764e-39 = -1.42174e-38
	(b"00000000011110010011111110110011", b"00000000000000000000000000000000"),
	(b"00000000001000111110111001101100", b"00000000100111010010111000011111"), -- 1.11349e-38 + 3.29977e-39 = 1.44347e-38
	(b"00000000000110001111001011111010", b"00000000000000000000000000000000"),
	(b"10000000001001001010001000100100", b"10000000000010111010111100101010"), -- 2.29122e-39 + -3.36424e-39 = -1.07303e-39
	(b"10000000011110010001111001000011", b"00000000000000000000000000000000"),
	(b"10000000010011101000100010110110", b"10000000110001111010011011111001"), -- -1.1123e-38 + -7.21221e-39 = -1.83352e-38
	(b"10000000001001111101001101010100", b"00000000000000000000000000000000"),
	(b"00000000000010100101101011100101", b"10000000000111010111100001101111"), -- -3.65739e-39 + 9.50962e-40 = -2.70643e-39
	(b"00000000001100011010010001000101", b"00000000000000000000000000000000"),
	(b"00000000001001000100101011000001", b"00000000010101011110111100000110"), -- 4.55887e-39 + 3.33289e-39 = 7.89176e-39
	(b"00000000001101011010101101011011", b"00000000000000000000000000000000"),
	(b"10000000001000100101110001011111", b"00000000000100110100111011111100"), -- 4.92875e-39 + -3.15554e-39 = 1.77321e-39
	(b"00000000001000011100111110000101", b"00000000000000000000000000000000"),
	(b"00000000001001000011110100111000", b"00000000010001100000110010111101"), -- 3.10502e-39 + 3.32804e-39 = 6.43305e-39
	(b"00000000010110011001100101011001", b"00000000000000000000000000000000"),
	(b"00000000000010111101111100111100", b"00000000011001010111100010010101"), -- 8.22837e-39 + 1.09027e-39 = 9.31864e-39
	(b"10000000001011001101111000001110", b"00000000000000000000000000000000"),
	(b"10000000011110101010101111010001", b"10000000101001111000100111011111"), -- -4.12042e-39 + -1.12656e-38 = -1.5386e-38
	(b"00000000001011011100111101011001", b"00000000000000000000000000000000"),
	(b"10000000001110000010110101001010", b"10000000000010100101110111110001"), -- 4.20698e-39 + -5.15903e-39 = -9.52055e-40
	(b"00000000001000010100111100111110", b"00000000000000000000000000000000"),
	(b"10000000001001000100011111111000", b"10000000000000101111100010111010"), -- 3.059e-39 + -3.3319e-39 = -2.72897e-40
	(b"00000000011010110111010011010101", b"00000000000000000000000000000000"),
	(b"10000000011100110111001110110100", b"10000000000001111111111011011111"), -- 9.86831e-39 + -1.06026e-38 = -7.34279e-40
	(b"00000000001100101101001100110100", b"00000000000000000000000000000000"),
	(b"10000000011111111001011101110001", b"10000000010011001100010000111101"), -- 4.66754e-39 + -1.17174e-38 = -7.04989e-39
	(b"10000000010101110110001110101001", b"00000000000000000000000000000000"),
	(b"10000000000101100011010010001101", b"10000000011011011001100000110110"), -- -8.02544e-39 + -2.03923e-39 = -1.00647e-38
	(b"10000000001110001000100000010001", b"00000000000000000000000000000000"),
	(b"00000000001000010111100001001110", b"10000000000101110000111111000011"), -- -5.1916e-39 + 3.07373e-39 = -2.11787e-39
	(b"10000000010010101100010010000110", b"00000000000000000000000000000000"),
	(b"10000000010110100000011011010010", b"10000000101001001100101101011000"), -- -6.86633e-39 + -8.26764e-39 = -1.5134e-38
	(b"00000000000001110000000010101100", b"00000000000000000000000000000000"),
	(b"00000000001110110100011101111110", b"00000000010000100100100000101010"), -- 6.43089e-40 + 5.44394e-39 = 6.08703e-39
	(b"10000000000101001111111010011000", b"00000000000000000000000000000000"),
	(b"00000000010010000001011011101111", b"00000000001100110001100001010111"), -- -1.92804e-39 + 6.62038e-39 = 4.69234e-39
	(b"00000000011001111000000011000111", b"00000000000000000000000000000000"),
	(b"00000000011110100011001010110110", b"00000000111000011011001101111101"), -- 9.50525e-39 + 1.12221e-38 = 2.07274e-38
	(b"00000000001111101010101000111101", b"00000000000000000000000000000000"),
	(b"00000000001010111000101100100001", b"00000000011010100011010101011110"), -- 5.75487e-39 + 3.99884e-39 = 9.75371e-39
	(b"00000000011111001110111011101010", b"00000000000000000000000000000000"),
	(b"00000000010111010011010001010111", b"00000000110110100010001101000001"), -- 1.14733e-38 + 8.55948e-39 = 2.00328e-38
	(b"00000000001010111010011101000111", b"00000000000000000000000000000000"),
	(b"10000000011001111110010100111011", b"10000000001111000011110111110100"), -- 4.00893e-39 + -9.54129e-39 = -5.53235e-39
	(b"00000000000000101000101111001111", b"00000000000000000000000000000000"),
	(b"10000000011110011010010101001111", b"10000000011101110001100110000000"), -- 2.33825e-40 + -1.11714e-38 = -1.09376e-38
	(b"00000000000000101101000101010101", b"00000000000000000000000000000000"),
	(b"00000000011011001010101101101010", b"00000000011011110111110010111111"), -- 2.58765e-40 + 9.97973e-39 = 1.02385e-38
	(b"00000000000111110000001110010000", b"00000000000000000000000000000000"),
	(b"00000000001101011011011010111011", b"00000000010101001011101001001011"), -- 2.84818e-39 + 4.93283e-39 = 7.78101e-39
	(b"00000000010001101010110101000110", b"00000000000000000000000000000000"),
	(b"00000000010111100001001111111111", b"00000000101001001100000101000101"), -- 6.49064e-39 + 8.63971e-39 = 1.51304e-38
	(b"10000000011111100010001101111110", b"00000000000000000000000000000000"),
	(b"00000000000101001011001101000000", b"10000000011010010111000000111110"), -- -1.1584e-38 + 1.90101e-39 = -9.68299e-39
	(b"00000000000011110000100101011110", b"00000000000000000000000000000000"),
	(b"00000000011001010110010101001110", b"00000000011101000110111010101100"), -- 1.38089e-39 + 9.31173e-39 = 1.06926e-38
	(b"00000000001010001000011101011000", b"00000000000000000000000000000000"),
	(b"10000000001001101110011110110111", b"00000000000000011001111110100001"), -- 3.72197e-39 + -3.57287e-39 = 1.491e-40
	(b"00000000001011001010011100100100", b"00000000000000000000000000000000"),
	(b"00000000011001111010010101100010", b"00000000100101000100110010000110"), -- 4.10072e-39 + 9.51838e-39 = 1.36191e-38
	(b"10000000010011100110111001000000", b"00000000000000000000000000000000"),
	(b"00000000011111010010100101010111", b"00000000001011101011101100010111"), -- -7.20272e-39 + 1.14943e-38 = 4.29155e-39
	(b"00000000001101110100011011011100", b"00000000000000000000000000000000"),
	(b"10000000001101101000101001011101", b"00000000000000001011110001111111"), -- 5.07637e-39 + -5.00875e-39 = 6.76197e-41
	(b"10000000001011010001110100110100", b"00000000000000000000000000000000"),
	(b"10000000010101000001101100111110", b"10000000100000010011100001110010"), -- -4.14307e-39 + -7.72395e-39 = -1.1867e-38
	(b"10000000011100001010101101010111", b"00000000000000000000000000000000"),
	(b"10000000011011101110101110110101", b"10000000110111111001011100001100"), -- -1.0347e-38 + -1.01865e-38 = -2.05335e-38
	(b"10000000001000011100011010010111", b"00000000000000000000000000000000"),
	(b"00000000011011000001111010110001", b"00000000010010100101100000011010"), -- -3.10181e-39 + 9.92924e-39 = 6.82743e-39
	(b"10000000010110011010110111010000", b"00000000000000000000000000000000"),
	(b"00000000010010001010010111010101", b"10000000000100010000011111111011"), -- -8.23571e-39 + 6.67165e-39 = -1.56407e-39
	(b"10000000011101001100001011100010", b"00000000000000000000000000000000"),
	(b"00000000010101100100100011100001", b"10000000000111100111101000000001"), -- -1.07228e-38 + 7.924e-39 = -2.79883e-39
	(b"10000000011101111110011010100011", b"00000000000000000000000000000000"),
	(b"10000000000101001100000001001000", b"10000000100011001010011011101011"), -- -1.10112e-38 + -1.90569e-39 = -1.29168e-38
	(b"00000000001100101111110010101011", b"00000000000000000000000000000000"),
	(b"00000000001110111100110011100101", b"00000000011011101100100110010000"), -- 4.68241e-39 + 5.4918e-39 = 1.01742e-38
	(b"00000000011110110010101011110101", b"00000000000000000000000000000000"),
	(b"10000000010010111001100001010010", b"00000000001011111001001010100011"), -- 1.13112e-38 + -6.9423e-39 = 4.36887e-39
	(b"00000000000011011110001011100101", b"00000000000000000000000000000000"),
	(b"00000000010010000110110000110101", b"00000000010101100100111100011010"), -- 1.27526e-39 + 6.65097e-39 = 7.92623e-39
	(b"10000000010111000100010001000100", b"00000000000000000000000000000000"),
	(b"00000000010111010000111001100101", b"00000000000000001100101000100001"), -- -8.47335e-39 + 8.54586e-39 = 7.25102e-41
	(b"00000000011010110110100010000010", b"00000000000000000000000000000000"),
	(b"00000000000000111010100000111100", b"00000000011011110001000010111110"), -- 9.86389e-39 + 3.35858e-40 = 1.01997e-38
	(b"10000000000111111000111111100010", b"00000000000000000000000000000000"),
	(b"00000000011010101001111101111100", b"00000000010010110000111110011010"), -- -2.89852e-39 + 9.79177e-39 = 6.89326e-39
	(b"10000000001010011001001110111010", b"00000000000000000000000000000000"),
	(b"00000000000011010001010111000010", b"10000000000111000111110111111000"), -- -3.81825e-39 + 1.20167e-39 = -2.61658e-39
	(b"10000000010101101111000110100111", b"00000000000000000000000000000000"),
	(b"00000000011101011111011100011100", b"00000000000111110000010101110101"), -- -7.98454e-39 + 1.08334e-38 = 2.84886e-39
	(b"10000000000001011101101101001011", b"00000000000000000000000000000000"),
	(b"00000000001100111101100001000001", b"00000000001011011111110011110110"), -- -5.37845e-40 + 4.76119e-39 = 4.22334e-39
	(b"00000000010010101001111011100011", b"00000000000000000000000000000000"),
	(b"00000000001110000000111111111111", b"00000000100000101010111011100010"), -- 6.85282e-39 + 5.14853e-39 = 1.20014e-38
	(b"10000000001011010110101110100000", b"00000000000000000000000000000000"),
	(b"00000000001110110111011011001111", b"00000000000011100000101100101111"), -- -4.17121e-39 + 5.46091e-39 = 1.28971e-39
	(b"10000000000010011010101010011011", b"00000000000000000000000000000000"),
	(b"00000000011110100111101101001111", b"00000000011100001101000010110100"), -- -8.87721e-40 + 1.12482e-38 = 1.03604e-38
	(b"10000000011000100000111000110110", b"00000000000000000000000000000000"),
	(b"00000000010011100100001011100100", b"10000000000100111100101101010010"), -- -9.00498e-39 + 7.18716e-39 = -1.81781e-39
	(b"00000000010100111010111011101110", b"00000000000000000000000000000000"),
	(b"00000000000011011110000101101000", b"00000000011000011001000001010110"), -- 7.6851e-39 + 1.27472e-39 = 8.95982e-39
	(b"10000000011111111111101100001000", b"00000000000000000000000000000000"),
	(b"10000000001010001001001100000001", b"10000000101010001000111000001001"), -- -1.17532e-38 + -3.72615e-39 = -1.54793e-38
	(b"10000000011001110000110010100110", b"00000000000000000000000000000000"),
	(b"10000000001001000111110110000100", b"10000000100010111000101000101010"), -- -9.46359e-39 + -3.3511e-39 = -1.28147e-38
	(b"00000000010111000100001110001100", b"00000000000000000000000000000000"),
	(b"10000000000011011100010111000000", b"00000000010011100111110111001100"), -- 8.4731e-39 + -1.2648e-39 = 7.2083e-39
	(b"10000000010111011100010000010001", b"00000000000000000000000000000000"),
	(b"10000000001110110101010000101110", b"10000000100110010001100000111111"), -- -8.61104e-39 + -5.44849e-39 = -1.40595e-38
	(b"00000000001001110101001011110101", b"00000000000000000000000000000000"),
	(b"10000000000100100111011001111110", b"00000000000101001101110001110111"), -- 3.61134e-39 + -1.69555e-39 = 1.9158e-39
	(b"10000000010110001000100110101010", b"00000000000000000000000000000000"),
	(b"00000000010101100011010010111010", b"10000000000000100101010011110000"), -- -8.13091e-39 + 7.91677e-39 = -2.14141e-40
	(b"00000000011101001001111100011110", b"00000000000000000000000000000000"),
	(b"00000000000110100100010000110000", b"00000000100011101110001101001110"), -- 1.071e-38 + 2.41218e-39 = 1.31222e-38
	(b"10000000010100011110111001011101", b"00000000000000000000000000000000"),
	(b"00000000000001000100000110001011", b"10000000010011011010110011010010"), -- -7.52418e-39 + 3.90854e-40 = -7.13333e-39
	(b"10000000011001110000010011110111", b"00000000000000000000000000000000"),
	(b"10000000011001001100011100000111", b"10000000110010111100101111111110"), -- -9.46084e-39 + -9.25495e-39 = -1.87158e-38
	(b"10000000011110110111100011000100", b"00000000000000000000000000000000"),
	(b"00000000010010011000111111100010", b"10000000001100011110100011100010"), -- -1.13391e-38 + 6.75561e-39 = -4.58348e-39
	(b"00000000000100010011110100100110", b"00000000000000000000000000000000"),
	(b"10000000011001000011000011000000", b"10000000010100101111001110011010"), -- 1.58314e-39 + -9.20104e-39 = -7.6179e-39
	(b"10000000001011101001010111000101", b"00000000000000000000000000000000"),
	(b"00000000011110011111001110110010", b"00000000010010110101110111101101"), -- -4.27816e-39 + 1.11995e-38 = 6.92136e-39
	(b"00000000010011011011111001001000", b"00000000000000000000000000000000"),
	(b"10000000010110001111000101010011", b"10000000000010110011001100001011"), -- 7.13959e-39 + -8.16809e-39 = -1.0285e-39
	(b"10000000011101101010001101110101", b"00000000000000000000000000000000"),
	(b"10000000001011111011101111000011", b"10000000101001100101111100111000"), -- -1.08952e-38 + -4.38362e-39 = -1.52789e-38
	(b"00000000001000001110100100001000", b"00000000000000000000000000000000"),
	(b"10000000010100110101101011001111", b"10000000001100100111000111000111"), -- 3.02233e-39 + -7.65492e-39 = -4.63259e-39
	(b"10000000000101110111111001111011", b"00000000000000000000000000000000"),
	(b"00000000001011100100011100010010", b"00000000000101101100100010010111"), -- -2.15759e-39 + 4.24993e-39 = 2.09234e-39
	(b"10000000001100100101010000010111", b"00000000000000000000000000000000"),
	(b"10000000000001111111001111000111", b"10000000001110100100011111011110"), -- -4.62194e-39 + -7.30299e-40 = -5.35224e-39
	(b"00000000010000010010000110011011", b"00000000000000000000000000000000"),
	(b"00000000010001010001110111010011", b"00000000100001100011111101101110"), -- 5.98136e-39 + 6.34735e-39 = 1.23287e-38
	(b"00000000011111100011011011101110", b"00000000000000000000000000000000"),
	(b"10000000011110000011000110101011", b"00000000000001100000010101000011"), -- 1.1591e-38 + -1.10381e-38 = 5.52901e-40
	(b"00000000010000001011101011000111", b"00000000000000000000000000000000"),
	(b"00000000000011111110100001001001", b"00000000010100001010001100010000"), -- 5.94447e-39 + 1.46086e-39 = 7.40534e-39
	(b"10000000001101001011110001001010", b"00000000000000000000000000000000"),
	(b"10000000010110111110011101110010", b"10000000100100001010001110111100"), -- -4.84299e-39 + -8.44006e-39 = -1.3283e-38
	(b"00000000011101001001111111111001", b"00000000000000000000000000000000"),
	(b"10000000000100101011011000100001", b"00000000011000011110100111011000"), -- 1.07103e-38 + -1.71837e-39 = 8.99193e-39
	(b"10000000001101000010110101110111", b"00000000000000000000000000000000"),
	(b"10000000010101111001010001100111", b"10000000100010111100000111011110"), -- -4.79176e-39 + -8.04292e-39 = -1.28347e-38
	(b"10000000011001001001001001100100", b"00000000000000000000000000000000"),
	(b"00000000010010111001001110100111", b"10000000000110001111111010111101"), -- -9.23606e-39 + 6.94063e-39 = -2.29543e-39
	(b"10000000011110001011001000010110", b"00000000000000000000000000000000"),
	(b"10000000010010100101011110010100", b"10000000110000110000100110101010"), -- -1.10841e-38 + -6.82724e-39 = -1.79114e-38
	(b"10000000000110000101001000101010", b"00000000000000000000000000000000"),
	(b"10000000011100010100000110111100", b"10000000100010011001001111100110"), -- -2.23353e-39 + -1.0401e-38 = -1.26345e-38
	(b"00000000011110101011111000110110", b"00000000000000000000000000000000"),
	(b"00000000000100001111100010011001", b"00000000100010111011011011001111"), -- 1.12722e-38 + 1.55855e-39 = 1.28307e-38
	(b"00000000001010100000110111100000", b"00000000000000000000000000000000"),
	(b"00000000000000111111011101101010", b"00000000001011100000010101001010"), -- 3.86207e-39 + 3.64262e-40 = 4.22633e-39
	(b"00000000000111001011111001110011", b"00000000000000000000000000000000"),
	(b"00000000000000001001010001010111", b"00000000000111010101001011001010"), -- 2.63971e-39 + 5.32143e-41 = 2.69293e-39
	(b"00000000000111110101000111000011", b"00000000000000000000000000000000"),
	(b"10000000011111100001000011110110", b"10000000010111101011111100110011"), -- 2.87623e-39 + -1.15774e-38 = -8.70113e-39
	(b"10000000010000101101010010111100", b"00000000000000000000000000000000"),
	(b"10000000001001101110100100100011", b"10000000011010011011110111011111"), -- -6.13746e-39 + -3.57338e-39 = -9.71084e-39
	(b"10000000011100011010000000110100", b"00000000000000000000000000000000"),
	(b"00000000011101011100011101001101", b"00000000000001000010011100011001"), -- -1.04349e-38 + 1.08162e-38 = 3.81368e-40
	(b"10000000011010001010010110011010", b"00000000000000000000000000000000"),
	(b"00000000000000000101000000000101", b"10000000011010000101010110010101"), -- -9.6103e-39 + 2.87056e-41 = -9.58159e-39
	(b"00000000011010001100101001000111", b"00000000000000000000000000000000"),
	(b"00000000000010010101111011000001", b"00000000011100100010100100001000"), -- 9.62346e-39 + 8.60511e-40 = 1.0484e-38
	(b"00000000000000100101110101010101", b"00000000000000000000000000000000"),
	(b"00000000011001101100011111001000", b"00000000011010010010010100011101"), -- 2.17152e-40 + 9.43889e-39 = 9.65604e-39
	(b"10000000010110110111101111011010", b"00000000000000000000000000000000"),
	(b"10000000001111100110111011011101", b"10000000100110011110101010110111"), -- -8.40146e-39 + -5.73357e-39 = -1.4135e-38
	(b"10000000011101000001000011000011", b"00000000000000000000000000000000"),
	(b"00000000000100111111000111101010", b"10000000011000000001111011011001"), -- -1.06589e-38 + 1.83166e-39 = -8.82727e-39
	(b"10000000011010101110000010101111", b"00000000000000000000000000000000"),
	(b"10000000010100101101010011101100", b"10000000101111011011010110011011"), -- -9.81516e-39 + -7.60689e-39 = -1.74221e-38
	(b"10000000011001100010110111101110", b"00000000000000000000000000000000"),
	(b"00000000011110111011100001000110", b"00000000000101011000101001011000"), -- -9.3837e-39 + 1.13619e-38 = 1.97817e-39
	(b"10000000001011010110100111111111", b"00000000000000000000000000000000"),
	(b"00000000011110000100011100001100", b"00000000010010101101110100001101"), -- -4.17062e-39 + 1.10457e-38 = 6.87512e-39
	(b"00000000010100011010100100111110", b"00000000000000000000000000000000"),
	(b"00000000010100000111001000010100", b"00000000101000100001101101010010"), -- 7.49939e-39 + 7.38776e-39 = 1.48872e-38
	(b"00000000000111101110101101101111", b"00000000000000000000000000000000"),
	(b"10000000001011111101000001001101", b"10000000000100001110010011011110"), -- 2.83952e-39 + -4.39099e-39 = -1.55147e-39
	(b"00000000011011100000001111101111", b"00000000000000000000000000000000"),
	(b"00000000010011100101001000001010", b"00000000101111000101010111111001"), -- 1.01033e-38 + 7.1926e-39 = 1.72959e-38
	(b"10000000010000101110101111010001", b"00000000000000000000000000000000"),
	(b"00000000001100010101110001110101", b"10000000000100011000111101011100"), -- -6.14574e-39 + 4.53311e-39 = -1.61263e-39
	(b"10000000001100100011101011100011", b"00000000000000000000000000000000"),
	(b"10000000000000100011000101101001", b"10000000001101000110110001001100"), -- -4.6129e-39 + -2.01396e-40 = -4.8143e-39
	(b"00000000011111110110001110111100", b"00000000000000000000000000000000"),
	(b"10000000010111101110100010110011", b"00000000001000000111101100001001"), -- 1.16989e-38 + -8.71601e-39 = 2.98287e-39
	(b"00000000000001101000110001000101", b"00000000000000000000000000000000"),
	(b"00000000000001001101011000100101", b"00000000000010110110001001101010"), -- 6.01332e-40 + 4.44163e-40 = 1.04549e-39
	(b"00000000011000101000110110011001", b"00000000000000000000000000000000"),
	(b"10000000001110011111110001101110", b"00000000001010001001000100101011"), -- 9.05067e-39 + -5.32518e-39 = 3.7255e-39
	(b"10000000011110011110010000010100", b"00000000000000000000000000000000"),
	(b"10000000000000000101110110101001", b"10000000011110100100000110111101"), -- -1.11939e-38 + -3.35989e-41 = -1.12275e-38
	(b"10000000001100110111010101100111", b"00000000000000000000000000000000"),
	(b"10000000001011010100001000010100", b"10000000011000001011011101111011"), -- -4.72573e-39 + -4.1563e-39 = -8.88203e-39
	(b"10000000010100100010010111000111", b"00000000000000000000000000000000"),
	(b"10000000001111011000001011001101", b"10000000100011111010100010010100"), -- -7.54406e-39 + -5.64889e-39 = -1.3193e-38
	(b"00000000010101100010101010011010", b"00000000000000000000000000000000"),
	(b"00000000000111001011010001111011", b"00000000011100101101111100010101"), -- 7.91314e-39 + 2.63614e-39 = 1.05493e-38
	(b"10000000011010111111110011100001", b"00000000000000000000000000000000"),
	(b"00000000000101010100111101111011", b"10000000010101101010110101100110"), -- -9.91711e-39 + 1.95706e-39 = -7.96006e-39
	(b"10000000011000100011101100110111", b"00000000000000000000000000000000"),
	(b"00000000001110101100010010011000", b"10000000001001110111011010011111"), -- -9.02112e-39 + 5.39698e-39 = -3.62414e-39
	(b"10000000011110011100110010011110", b"00000000000000000000000000000000"),
	(b"10000000001010010101100000000111", b"10000000101000110010010010100101"), -- -1.11855e-38 + -3.79683e-39 = -1.49823e-38
	(b"10000000000011001010000011101100", b"00000000000000000000000000000000"),
	(b"00000000011100000010110011010101", b"00000000011000111000101111101001"), -- -1.15975e-39 + 1.03017e-38 = 9.1419e-39
	(b"10000000011001101100000010110011", b"00000000000000000000000000000000"),
	(b"10000000000010101001100011011110", b"10000000011100010101100110010001"), -- -9.43635e-39 + -9.73193e-40 = -1.04095e-38
	(b"10000000001011111000011100000001", b"00000000000000000000000000000000"),
	(b"10000000001011011100110010100101", b"10000000010111010101001110100110"), -- -4.3647e-39 + -4.20601e-39 = -8.57071e-39
	(b"10000000000101010011010100101100", b"00000000000000000000000000000000"),
	(b"10000000010101110100011011111110", b"10000000011011000111110000101010"), -- -1.94762e-39 + -8.01516e-39 = -9.96278e-39
	(b"00000000001011111011000011001010", b"00000000000000000000000000000000"),
	(b"10000000011100010110111111110001", b"10000000010000011011111100100111"), -- 4.37969e-39 + -1.04176e-38 = -6.03788e-39
	(b"10000000010011111010100101100100", b"00000000000000000000000000000000"),
	(b"10000000000100110100100101011110", b"10000000011000101111001011000010"), -- -7.31577e-39 + -1.77119e-39 = -9.08696e-39
	(b"00000000000001110100100010010101", b"00000000000000000000000000000000"),
	(b"00000000010011101001111010111111", b"00000000010101011110011101010100"), -- 6.68886e-40 + 7.22012e-39 = 7.889e-39
	(b"10000000010100000111100101011101", b"00000000000000000000000000000000"),
	(b"10000000001110011001010000000010", b"10000000100010100000110101011111"), -- -7.39038e-39 + -5.28772e-39 = -1.26781e-38
	(b"10000000001000000000001001000010", b"00000000000000000000000000000000"),
	(b"10000000000101110000001100111010", b"10000000001101110000010101111100"), -- -2.93955e-39 + -2.11337e-39 = -5.05292e-39
	(b"10000000011001101001110101010010", b"00000000000000000000000000000000"),
	(b"10000000001110101111101101011010", b"10000000101000011001100010101100"), -- -9.42366e-39 + -5.41663e-39 = -1.48403e-38
	(b"00000000011100110111101101000000", b"00000000000000000000000000000000"),
	(b"00000000001110000001001001110101", b"00000000101010111000110110110101"), -- 1.06053e-38 + 5.14941e-39 = 1.57547e-38
	(b"00000000000011100110000111100101", b"00000000000000000000000000000000"),
	(b"10000000001010100101000010011000", b"10000000000110111110111010110011"), -- 1.32081e-39 + -3.886e-39 = -2.56519e-39
	(b"10000000011101110000101101000100", b"00000000000000000000000000000000"),
	(b"10000000001110010011010011110111", b"10000000101100000100000000111011"), -- -1.09325e-38 + -5.25362e-39 = -1.61861e-38
	(b"00000000011001111000000101010011", b"00000000000000000000000000000000"),
	(b"10000000001001111001001011001100", b"00000000001111111110111010000111"), -- 9.50545e-39 + -3.63425e-39 = 5.8712e-39
	(b"10000000011000110001110100101101", b"00000000000000000000000000000000"),
	(b"10000000000100000100011110000011", b"10000000011100110110010010110000"), -- -9.10218e-39 + -1.49502e-39 = -1.05972e-38
	(b"00000000010101011000110011101111", b"00000000000000000000000000000000"),
	(b"10000000000100000010001000101101", b"00000000010001010110101011000010"), -- 7.85657e-39 + -1.48163e-39 = 6.37495e-39
	(b"10000000000110010001011100010100", b"00000000000000000000000000000000"),
	(b"10000000010101011100010010101101", b"10000000011011101101101111000001"), -- -2.30417e-39 + -7.87657e-39 = -1.01807e-38
	(b"10000000001110011100100000010110", b"00000000000000000000000000000000"),
	(b"00000000001000100101000000110011", b"10000000000101110111011111100011"), -- -5.3064e-39 + 3.15118e-39 = -2.15522e-39
	(b"00000000011101001001101001110010", b"00000000000000000000000000000000"),
	(b"00000000011011000000001111010001", b"00000000111000001001111001000011"), -- 1.07083e-38 + 9.9196e-39 = 2.06279e-38
	(b"10000000001111101010101110001101", b"00000000000000000000000000000000"),
	(b"00000000000111110111011010000011", b"10000000000111110011010100001010"), -- -5.75534e-39 + 2.88941e-39 = -2.86593e-39
	(b"00000000010000100010110001010111", b"00000000000000000000000000000000"),
	(b"00000000000010001001110111110001", b"00000000010010101100101001001000"), -- 6.07705e-39 + 7.91343e-40 = 6.86839e-39
	(b"10000000010010011001011011011100", b"00000000000000000000000000000000"),
	(b"00000000010010011111010110101010", b"00000000000000000101111011001110"), -- -6.75811e-39 + 6.79212e-39 = 3.40095e-41
	(b"10000000010110000110100000100110", b"00000000000000000000000000000000"),
	(b"10000000000001000101010000110001", b"10000000010111001011110001010111"), -- -8.11889e-39 + -3.97544e-40 = -8.51643e-39
	(b"00000000001001100010010001011011", b"00000000000000000000000000000000"),
	(b"10000000000100110000010010000000", b"00000000000100110001111111011011"), -- 3.50279e-39 + -1.74649e-39 = 1.7563e-39
	(b"00000000001001010110100111010101", b"00000000000000000000000000000000"),
	(b"10000000010000010010110110001010", b"10000000000110111100001110110101"), -- 3.43588e-39 + -5.98564e-39 = -2.54976e-39
	(b"10000000001111011000110110111110", b"00000000000000000000000000000000"),
	(b"10000000010110101000010101010000", b"10000000100110000001001100001110"), -- -5.65281e-39 + -8.31302e-39 = -1.39658e-38
	(b"00000000000101010111110101010011", b"00000000000000000000000000000000"),
	(b"00000000011011100110111010110101", b"00000000100000111110110000001000"), -- 1.9735e-39 + 1.01416e-38 = 1.21151e-38
	(b"00000000010101001001010011110100", b"00000000000000000000000000000000"),
	(b"10000000011101000100101010110000", b"10000000000111111011010110111100"), -- 7.76762e-39 + -1.06797e-38 = -2.91209e-39
	(b"00000000011010010110011001110011", b"00000000000000000000000000000000"),
	(b"10000000000000010110111011101110", b"00000000011001111111011110000101"), -- 9.67948e-39 + -1.3163e-40 = 9.54785e-39
	(b"10000000001001001111010100101000", b"00000000000000000000000000000000"),
	(b"10000000010111100100000000010100", b"10000000100000110011010100111100"), -- -3.39402e-39 + -8.65552e-39 = -1.20495e-38
	(b"00000000010000011101100000101100", b"00000000000000000000000000000000"),
	(b"10000000011100110011101001010101", b"10000000001100010110001000101001"), -- 6.04686e-39 + -1.0582e-38 = -4.53515e-39
	(b"10000000000111111101011100000110", b"00000000000000000000000000000000"),
	(b"00000000011110000000000010100001", b"00000000010110000010100110011011"), -- -2.92404e-39 + 1.10205e-38 = 8.09645e-39
	(b"00000000010110111110110010101111", b"00000000000000000000000000000000"),
	(b"00000000011011100110110000101101", b"00000000110010100101100011011100"), -- 8.44194e-39 + 1.01407e-38 = 1.85826e-38
	(b"00000000010011111110000011111111", b"00000000000000000000000000000000"),
	(b"00000000000001011010011100100001", b"00000000010101011000100000100000"), -- 7.33572e-39 + 5.19132e-40 = 7.85485e-39
	(b"10000000011101010010110011000101", b"00000000000000000000000000000000"),
	(b"00000000000110111010000001011101", b"10000000010110011000110001101000"), -- -1.07608e-38 + 2.53709e-39 = -8.22373e-39
	(b"10000000000000010111000110110101", b"00000000000000000000000000000000"),
	(b"00000000011001110101110010101001", b"00000000011001011110101011110100"), -- -1.32626e-40 + 9.4923e-39 = 9.35967e-39
	(b"00000000010101110001101101001101", b"00000000000000000000000000000000"),
	(b"10000000000011010010001000010010", b"00000000010010011111100100111011"), -- 7.99948e-39 + -1.20608e-39 = 6.7934e-39
	(b"00000000011011101100010101001010", b"00000000000000000000000000000000"),
	(b"10000000010011111001100001001000", b"00000000000111110010110100000010"), -- 1.01727e-38 + -7.30963e-39 = 2.86305e-39
	(b"10000000000111011010101110110101", b"00000000000000000000000000000000"),
	(b"00000000001011001000011111101101", b"00000000000011101101110000111000"), -- -2.72483e-39 + 4.08952e-39 = 1.3647e-39
	(b"10000000010011011101001010110010", b"00000000000000000000000000000000"),
	(b"00000000010011011100100110001001", b"10000000000000000000100100101001"), -- -7.14692e-39 + 7.14363e-39 = -3.28604e-42
	(b"10000000010110001011100011000110", b"00000000000000000000000000000000"),
	(b"10000000000011010000011100100101", b"10000000011001011011111111101011"), -- -8.14781e-39 + -1.19642e-39 = -9.34423e-39
	(b"00000000001010011010010000000101", b"00000000000000000000000000000000"),
	(b"00000000000101100011011111111101", b"00000000001111111101110000000010"), -- 3.82409e-39 + 2.04047e-39 = 5.86456e-39
	(b"00000000001101100110000010100111", b"00000000000000000000000000000000"),
	(b"00000000001100000010100001000100", b"00000000011001101000100011101011"), -- 4.99379e-39 + 4.42255e-39 = 9.41634e-39
	(b"10000000011001010010100011001001", b"00000000000000000000000000000000"),
	(b"00000000011111011101101010001001", b"00000000000110001011000111000000"), -- -9.29002e-39 + 1.15578e-38 = 2.26782e-39
	(b"00000000011001001011000111101010", b"00000000000000000000000000000000"),
	(b"00000000000110111110111010010100", b"00000000100000001010000001111110"), -- 9.24737e-39 + 2.56514e-39 = 1.18125e-38
	(b"00000000010111000101111111110111", b"00000000000000000000000000000000"),
	(b"10000000010110101101010100011000", b"00000000000000011000101011011111"), -- 8.48329e-39 + -8.34164e-39 = 1.41653e-40
	(b"00000000010101110001101100001001", b"00000000000000000000000000000000"),
	(b"00000000010111100010010111101101", b"00000000101101010100000011110110"), -- 7.99939e-39 + 8.64614e-39 = 1.66455e-38
	(b"00000000000011000100010010111001", b"00000000000000000000000000000000"),
	(b"00000000011001100000001000111000", b"00000000011100100100011011110001"), -- 1.12668e-39 + 9.36802e-39 = 1.04947e-38
	(b"10000000000101100001011100110001", b"00000000000000000000000000000000"),
	(b"10000000010010100100000101111010", b"10000000011000000101100010101011"), -- -2.0287e-39 + -6.81932e-39 = -8.84802e-39
	(b"00000000000011000001010010110001", b"00000000000000000000000000000000"),
	(b"00000000010010101100001010101101", b"00000000010101101101011101011110"), -- 1.10945e-39 + 6.86566e-39 = 7.97511e-39
	(b"00000000000110101001000100111100", b"00000000000000000000000000000000"),
	(b"00000000000001110001110001011001", b"00000000001000011010110110010101"), -- 2.43982e-39 + 6.53018e-40 = 3.09284e-39
	(b"00000000011011010110001000001101", b"00000000000000000000000000000000"),
	(b"10000000001001000110111010100100", b"00000000010010001111001101101001"), -- 1.00452e-38 + -3.34577e-39 = 6.69947e-39
	(b"00000000000111111010001111000100", b"00000000000000000000000000000000"),
	(b"00000000001111111001100011010000", b"00000000010111110011110010010100"), -- 2.90565e-39 + 5.84046e-39 = 8.7461e-39
	(b"10000000000001001100111100001101", b"00000000000000000000000000000000"),
	(b"00000000001000000100100011010000", b"00000000000110110111100111000011"), -- -4.41618e-40 + 2.96486e-39 = 2.52324e-39
	(b"10000000001111010111000100011111", b"00000000000000000000000000000000"),
	(b"00000000000100111101101111001111", b"10000000001010011001010101010000"), -- -5.64255e-39 + 1.82373e-39 = -3.81882e-39
	(b"00000000010111010010111101110110", b"00000000000000000000000000000000"),
	(b"00000000010101111110000111011011", b"00000000101101010001000101010001"), -- 8.55773e-39 + 8.07071e-39 = 1.66284e-38
	(b"10000000000111101010110011110011", b"00000000000000000000000000000000"),
	(b"10000000001010000101111111001000", b"10000000010001110000110010111011"), -- -2.81711e-39 + -3.70778e-39 = -6.52489e-39
	(b"00000000010000000101011100000011", b"00000000000000000000000000000000"),
	(b"00000000001010110001111100011000", b"00000000011010110111011000011011"), -- 5.90869e-39 + 3.96008e-39 = 9.86877e-39
	(b"10000000001110010101010110000010", b"00000000000000000000000000000000"),
	(b"10000000001010111011111001111101", b"10000000011001010001001111111111"), -- -5.2653e-39 + -4.01726e-39 = -9.28256e-39
	(b"10000000000110010000011000100010", b"00000000000000000000000000000000"),
	(b"10000000000101111101010001001010", b"10000000001100001101101001101100"), -- -2.29809e-39 + -2.18837e-39 = -4.48646e-39
	(b"00000000011100011000000000011010", b"00000000000000000000000000000000"),
	(b"10000000011011101111001110101000", b"00000000000000101000110001110010"), -- 1.04234e-38 + -1.01893e-38 = 2.34053e-40
	(b"00000000000110111111000111110110", b"00000000000000000000000000000000"),
	(b"00000000000011001101111110000000", b"00000000001010001101000101110110"), -- 2.56636e-39 + 1.1822e-39 = 3.74856e-39
	(b"00000000001100110101010001010010", b"00000000000000000000000000000000"),
	(b"00000000000000001010000000101110", b"00000000001100111111010010000000"), -- 4.71386e-39 + 5.74616e-41 = 4.77132e-39
	(b"10000000001000111110001011110110", b"00000000000000000000000000000000"),
	(b"10000000000010000011011000100110", b"10000000001011000001100100011100"), -- -3.29566e-39 + -7.54109e-40 = -4.04977e-39
	(b"10000000000101111010111101101000", b"00000000000000000000000000000000"),
	(b"00000000010100000001100011111000", b"00000000001110000110100110010000"), -- -2.17514e-39 + 7.3558e-39 = 5.18066e-39
	(b"10000000001011001011011001100101", b"00000000000000000000000000000000"),
	(b"10000000000110011101000111001010", b"10000000010001101000100000101111"), -- -4.10619e-39 + -2.37115e-39 = -6.47734e-39
	(b"10000000011000101100111101101001", b"00000000000000000000000000000000"),
	(b"10000000001110000010011100000110", b"10000000100110101111011001101111"), -- -9.07428e-39 + -5.15679e-39 = -1.42311e-38
	(b"00000000001100000011101111110011", b"00000000000000000000000000000000"),
	(b"10000000010001111110001110001010", b"10000000000101111010011110010111"), -- 4.42961e-39 + -6.60195e-39 = -2.17234e-39
	(b"10000000001111101010101000111011", b"00000000000000000000000000000000"),
	(b"00000000010101001101001000000000", b"00000000000101100010011111000101"), -- -5.75487e-39 + 7.78952e-39 = 2.03465e-39
	(b"00000000010100100110101101000101", b"00000000000000000000000000000000"),
	(b"00000000010001010011110011110001", b"00000000100101111010100000110110"), -- 7.56899e-39 + 6.35851e-39 = 1.39275e-38
	(b"00000000010000010100111111100000", b"00000000000000000000000000000000"),
	(b"10000000001011001010100111010100", b"00000000000101001010011000001100"), -- 5.99796e-39 + -4.10168e-39 = 1.89628e-39
	(b"00000000010001101111100111101101", b"00000000000000000000000000000000"),
	(b"10000000001100000100111010001000", b"00000000000101101010101101100101"), -- 6.51814e-39 + -4.43628e-39 = 2.08187e-39
	(b"00000000000000111100111011000001", b"00000000000000000000000000000000"),
	(b"00000000010110000100101010100010", b"00000000010111000001100101100011"), -- 3.49676e-40 + 8.1083e-39 = 8.45797e-39
	(b"00000000001101001110101110010101", b"00000000000000000000000000000000"),
	(b"10000000011111111101010010110100", b"10000000010010101110100100011111"), -- 4.85996e-39 + -1.17394e-38 = -6.87945e-39
	(b"10000000001111111011000000010000", b"00000000000000000000000000000000"),
	(b"10000000000101110000101011110000", b"10000000010101101011101100000000"), -- -5.8488e-39 + -2.11614e-39 = -7.96494e-39
	(b"10000000010100011000001000110110", b"00000000000000000000000000000000"),
	(b"10000000000001101001011000110011", b"10000000010110000001100001101001"), -- -7.48539e-39 + -6.04894e-40 = -8.09028e-39
	(b"00000000011011010001010000100001", b"00000000000000000000000000000000"),
	(b"10000000001010111010111011011100", b"00000000010000010110010101000101"), -- 1.00173e-38 + -4.01165e-39 = 6.00564e-39
	(b"00000000010101000010101010011100", b"00000000000000000000000000000000"),
	(b"00000000001111100011110001010011", b"00000000100100100110011011101111"), -- 7.72947e-39 + 5.71544e-39 = 1.34449e-38
	(b"10000000011100101110011010010000", b"00000000000000000000000000000000"),
	(b"10000000010111001011101011111110", b"10000000110011111010000110001110"), -- -1.0552e-38 + -8.51595e-39 = -1.90679e-38
	(b"10000000011100010001001100111111", b"00000000000000000000000000000000"),
	(b"10000000011100011001111001100010", b"10000000111000101011000110100001"), -- -1.03843e-38 + -1.04342e-38 = -2.08185e-38
	(b"00000000000000110010001100100001", b"00000000000000000000000000000000"),
	(b"10000000011000111010100101000000", b"10000000011000001000011000011111"), -- 2.88108e-40 + -9.15243e-39 = -8.86432e-39
	(b"10000000010111010100011001011000", b"00000000000000000000000000000000"),
	(b"00000000011101111101111110100101", b"00000000000110101001100101001101"), -- -8.56594e-39 + 1.10087e-38 = 2.44272e-39
	(b"00000000000000010111001111011000", b"00000000000000000000000000000000"),
	(b"10000000011100001000101100011011", b"10000000011011110001011101000011"), -- 1.33392e-40 + -1.03355e-38 = -1.02021e-38
	(b"00000000011101011110011010110100", b"00000000000000000000000000000000"),
	(b"10000000000000111110100110101101", b"00000000011100011111110100000111"), -- 1.08275e-38 + -3.59334e-40 = 1.04682e-38
	(b"10000000001111011010111110111101", b"00000000000000000000000000000000"),
	(b"10000000011000101010101000110001", b"10000000101000000101100111101110"), -- -5.66501e-39 + -9.06093e-39 = -1.47259e-38
	(b"00000000011011011011100000011111", b"00000000000000000000000000000000"),
	(b"00000000011110101011100100100110", b"00000000111010000111000101000101"), -- 1.00761e-38 + 1.12703e-38 = 2.13465e-38
	(b"10000000010000111111110110010000", b"00000000000000000000000000000000"),
	(b"00000000010010011101101110010110", b"00000000000001011101111000000110"), -- -6.24394e-39 + 6.78276e-39 = 5.38824e-40
	(b"10000000011010101001100010101100", b"00000000000000000000000000000000"),
	(b"00000000011101101000001100110111", b"00000000000010111110101010001011"), -- -9.78933e-39 + 1.08837e-38 = 1.09433e-39
	(b"10000000000010100111011100111101", b"00000000000000000000000000000000"),
	(b"10000000001111001000000010011111", b"10000000010001101111011111011100"), -- -9.6113e-40 + -5.55627e-39 = -6.5174e-39
	(b"10000000001001100010101101000110", b"00000000000000000000000000000000"),
	(b"00000000000110111011001001110011", b"10000000000010100111100011010011"), -- -3.50527e-39 + 2.54357e-39 = -9.61699e-40
	(b"10000000001001001101110100010110", b"00000000000000000000000000000000"),
	(b"10000000011001000111001011101111", b"10000000100010010101000000000101"), -- -3.38539e-39 + -9.22478e-39 = -1.26102e-38
	(b"10000000000100011000101101101100", b"00000000000000000000000000000000"),
	(b"00000000010111000011010110000101", b"00000000010010101010101000011001"), -- -1.61122e-39 + 8.46806e-39 = 6.85685e-39
	(b"10000000001111101001100111011001", b"00000000000000000000000000000000"),
	(b"00000000001101010011001110000111", b"10000000000010010110011001010010"), -- -5.74899e-39 + 4.88577e-39 = -8.63225e-40
	(b"00000000010010101011000011100010", b"00000000000000000000000000000000"),
	(b"10000000000011111100111100111111", b"00000000001110101110000110100011"), -- 6.85928e-39 + -1.45188e-39 = 5.4074e-39
	(b"00000000000111011110000100110001", b"00000000000000000000000000000000"),
	(b"10000000010111110101001011111011", b"10000000010000010111000111001010"), -- 2.74401e-39 + -8.75414e-39 = -6.01013e-39
	(b"00000000010101111010110010100100", b"00000000000000000000000000000000"),
	(b"10000000000010011100001111110110", b"00000000010011011110100010101110"), -- 8.05162e-39 + -8.96817e-40 = 7.1548e-39
	(b"10000000011101011111111000100110", b"00000000000000000000000000000000"),
	(b"10000000011010101101000100001101", b"10000000111000001100111100110011"), -- -1.08359e-38 + -9.80956e-39 = -2.06455e-38
	(b"00000000010010100000011111110000", b"00000000000000000000000000000000"),
	(b"00000000000111100100001111011100", b"00000000011010000100101111001100"), -- 6.79867e-39 + 2.77941e-39 = 9.57808e-39
	(b"00000000001111011101010111100111", b"00000000000000000000000000000000"),
	(b"10000000010000000101110100111001", b"10000000000000101000011101010010"), -- 5.6787e-39 + -5.91091e-39 = -2.32215e-40
	(b"10000000011110001010000001001010", b"00000000000000000000000000000000"),
	(b"10000000011101101011001101011101", b"10000000111011110101001110100111"), -- -1.10778e-38 + -1.09009e-38 = -2.19787e-38
	(b"00000000000111110111110001111000", b"00000000000000000000000000000000"),
	(b"00000000001101000010011000000011", b"00000000010100111010001001111011"), -- 2.89155e-39 + 4.78908e-39 = 7.68063e-39
	(b"10000000010111100110100000011111", b"00000000000000000000000000000000"),
	(b"10000000010010011011000100010011", b"10000000101010000001100100110010"), -- -8.66989e-39 + -6.76751e-39 = -1.54374e-38
	(b"00000000001101100110111100111010", b"00000000000000000000000000000000"),
	(b"00000000000110011110101111101110", b"00000000010100000101101100101000"), -- 4.99902e-39 + 2.38052e-39 = 7.37954e-39
	(b"00000000011101110100101001111011", b"00000000000000000000000000000000"),
	(b"00000000010011111111101011010111", b"00000000110001110100010101010010"), -- 1.09551e-38 + 7.34499e-39 = 1.83001e-38
	(b"10000000010111001101101011110110", b"00000000000000000000000000000000"),
	(b"10000000000101011000011100010101", b"10000000011100100110001000001011"), -- -8.52741e-39 + -1.977e-39 = -1.05044e-38
	(b"00000000001010011010010000010010", b"00000000000000000000000000000000"),
	(b"10000000001111100100010101100111", b"10000000000101001010000101010101"), -- 3.82411e-39 + -5.7187e-39 = -1.89458e-39
	(b"00000000011101111000010101101000", b"00000000000000000000000000000000"),
	(b"10000000010111001111101111110100", b"00000000000110101000100101110100"), -- 1.09763e-38 + -8.53925e-39 = 2.43703e-39
	(b"10000000011100010010110110010110", b"00000000000000000000000000000000"),
	(b"10000000000101100010010000100110", b"10000000100001110101000110111100"), -- -1.03938e-38 + -2.03335e-39 = -1.24271e-38
	(b"10000000001101111011010101011110", b"00000000000000000000000000000000"),
	(b"10000000001111011010010110110111", b"10000000011101010101101100010101"), -- -5.11601e-39 + -5.66141e-39 = -1.07774e-38
	(b"10000000001110000100101010010110", b"00000000000000000000000000000000"),
	(b"00000000011001111101000001110010", b"00000000001011111000010111011100"), -- -5.16954e-39 + 9.53383e-39 = 4.36429e-39
	(b"10000000011110111010110011111101", b"00000000000000000000000000000000"),
	(b"00000000011010100010110010100010", b"10000000000100011000000001011011"), -- -1.13578e-38 + 9.75057e-39 = -1.60725e-39
	(b"10000000000001011000101001100111", b"00000000000000000000000000000000"),
	(b"00000000000000010011110000111110", b"10000000000001000100111000101001"), -- -5.08827e-40 + 1.13446e-40 = -3.95381e-40
	(b"00000000001001100100000010000100", b"00000000000000000000000000000000"),
	(b"00000000000101000011111010100110", b"00000000001110100111111100101010"), -- 3.51289e-39 + 1.85918e-39 = 5.37208e-39
	(b"10000000001000101011111100111110", b"00000000000000000000000000000000"),
	(b"10000000000110110111011100011001", b"10000000001111100011011001010111"), -- -3.19101e-39 + -2.52228e-39 = -5.71329e-39
	(b"00000000010001010010001100110110", b"00000000000000000000000000000000"),
	(b"00000000011110101010101111101101", b"00000000101111111100111100100011"), -- 6.34928e-39 + 1.12656e-38 = 1.76149e-38
	(b"00000000010100000101111110011110", b"00000000000000000000000000000000"),
	(b"00000000001001111011101111000010", b"00000000011110000001101101100000"), -- 7.38114e-39 + 3.64894e-39 = 1.10301e-38
	(b"10000000001000110101110110001011", b"00000000000000000000000000000000"),
	(b"00000000001111011110011011011000", b"00000000000110101000100101001101"), -- -3.2478e-39 + 5.68478e-39 = 2.43698e-39
	(b"00000000011111011111100011110010", b"00000000000000000000000000000000"),
	(b"00000000000110111100110101001010", b"00000000100110011100011000111100"), -- 1.15687e-38 + 2.5532e-39 = 1.41219e-38
	(b"00000000000011010000101010001001", b"00000000000000000000000000000000"),
	(b"00000000011100101000110010101100", b"00000000011111111001011100110101"), -- 1.19764e-39 + 1.05197e-38 = 1.17174e-38
	(b"10000000010010000101001000011101", b"00000000000000000000000000000000"),
	(b"00000000000010000111000100101001", b"10000000001111111110000011110100"), -- -6.64161e-39 + 7.75278e-40 = -5.86633e-39
	(b"10000000010110010001100000011111", b"00000000000000000000000000000000"),
	(b"00000000001000101001000101001100", b"10000000001101101000011011010011"), -- -8.18201e-39 + 3.17453e-39 = -5.00748e-39
	(b"00000000010011010111001000001001", b"00000000000000000000000000000000"),
	(b"10000000001100001000001010101100", b"00000000000111001110111101011101"), -- 7.11224e-39 + -4.45498e-39 = 2.65726e-39
	(b"10000000011001101000001010010110", b"00000000000000000000000000000000"),
	(b"00000000011101101101011101010100", b"00000000000100000101010010111110"), -- -9.41407e-39 + 1.09138e-38 = 1.49977e-39
	(b"00000000010001010100000110110111", b"00000000000000000000000000000000"),
	(b"00000000010100100101010001001101", b"00000000100101111001011000000100"), -- 6.36022e-39 + 7.56075e-39 = 1.3921e-38
	(b"10000000011010001011110011001001", b"00000000000000000000000000000000"),
	(b"00000000010000001000111111110111", b"10000000001010000010110011010010"), -- -9.61861e-39 + 5.92912e-39 = -3.6895e-39
	(b"10000000010111111111000110000011", b"00000000000000000000000000000000"),
	(b"10000000010110011100100100101100", b"10000000101110011011101010101111"), -- -8.81101e-39 + -8.24553e-39 = -1.70565e-38
	(b"10000000010011001110110001010011", b"00000000000000000000000000000000"),
	(b"10000000001010000101011001110010", b"10000000011101010100001011000101"), -- -7.06427e-39 + -3.70443e-39 = -1.07687e-38
	(b"00000000010111111011011011010111", b"00000000000000000000000000000000"),
	(b"00000000001001111001010110001010", b"00000000100001110100110001100001"), -- 8.78996e-39 + 3.63523e-39 = 1.24252e-38
	(b"00000000001011111101011000001111", b"00000000000000000000000000000000"),
	(b"00000000011110000110111001100101", b"00000000101010000100010001110100"), -- 4.39306e-39 + 1.10599e-38 = 1.54529e-38
	(b"00000000011001110001000111010111", b"00000000000000000000000000000000"),
	(b"00000000001101111011001101110111", b"00000000100111101100010101001110"), -- 9.46546e-39 + 5.11533e-39 = 1.45808e-38
	(b"10000000011101011100001110001001", b"00000000000000000000000000000000"),
	(b"10000000011111110100001111100101", b"10000000111101010000011101101110"), -- -1.08149e-38 + -1.16875e-38 = -2.25024e-38
	(b"00000000000011010001010101110110", b"00000000000000000000000000000000"),
	(b"00000000000010010011011111010110", b"00000000000101100100110101001100"), -- 1.20156e-39 + 8.4655e-40 = 2.04811e-39
	(b"00000000011011001001011011111111", b"00000000000000000000000000000000"),
	(b"10000000011111011111101011010000", b"10000000000100010110001111010001"), -- 9.9724e-39 + -1.15694e-38 = -1.59701e-39
	(b"00000000001011101011010001010111", b"00000000000000000000000000000000"),
	(b"00000000001010011101011111100010", b"00000000010110001000110000111001"), -- 4.28913e-39 + 3.8427e-39 = 8.13183e-39
	(b"00000000000110100111110111111000", b"00000000000000000000000000000000"),
	(b"10000000010110000000110111001111", b"10000000001111011000111111010111"), -- 2.43291e-39 + -8.08648e-39 = -5.65357e-39
	(b"00000000010010000011101011011010", b"00000000000000000000000000000000"),
	(b"00000000010010111100110001111111", b"00000000100101000000011101011001"), -- 6.63327e-39 + 6.96102e-39 = 1.35943e-38
	(b"00000000010010000111010101010100", b"00000000000000000000000000000000"),
	(b"10000000011010000111110111000101", b"10000000001000000000100001110001"), -- 6.65425e-39 + -9.59601e-39 = -2.94176e-39
	(b"10000000001101001101001010010111", b"00000000000000000000000000000000"),
	(b"00000000011010111100110100011011", b"00000000001101101111101010000100"), -- -4.85099e-39 + 9.89998e-39 = 5.04898e-39
	(b"00000000000001110100011111000101", b"00000000000000000000000000000000"),
	(b"00000000000100010010100000011110", b"00000000000110000110111111100011"), -- 6.68595e-40 + 1.57559e-39 = 2.24419e-39
	(b"00000000001001100000111111000111", b"00000000000000000000000000000000"),
	(b"10000000010010000101110110100111", b"10000000001000100100110111100000"), -- 3.49541e-39 + -6.64575e-39 = -3.15034e-39
	(b"10000000010000001111001001001011", b"00000000000000000000000000000000"),
	(b"10000000000111100101001001111011", b"10000000010111110100010011000110"), -- -5.96439e-39 + -2.78465e-39 = -8.74904e-39
	(b"10000000010111111001001100100011", b"00000000000000000000000000000000"),
	(b"10000000011011000011110100100100", b"10000000110010111101000001000111"), -- -8.77715e-39 + -9.94017e-39 = -1.87173e-38
	(b"10000000001111100111110100110001", b"00000000000000000000000000000000"),
	(b"00000000010110100100101110101011", b"00000000000110111100111001111010"), -- -5.73871e-39 + 8.29234e-39 = 2.55363e-39
	(b"00000000011100110100111100011100", b"00000000000000000000000000000000"),
	(b"10000000011100011100100111000101", b"00000000000000011000010101010111"), -- 1.05895e-38 + -1.04498e-38 = 1.39669e-40
	(b"00000000011110011011100110110010", b"00000000000000000000000000000000"),
	(b"00000000011011000000011100100110", b"00000000111001011100000011011000"), -- 1.11787e-38 + 9.9208e-39 = 2.10995e-38
	(b"10000000000111000001110111111110", b"00000000000000000000000000000000"),
	(b"00000000011000111001110101011011", b"00000000010001110111111101011101"), -- -2.58215e-39 + 9.14816e-39 = 6.56601e-39
	(b"10000000011011110010100110000111", b"00000000000000000000000000000000"),
	(b"00000000011111011000010011010011", b"00000000000011100101101101001100"), -- -1.02086e-38 + 1.15271e-38 = 1.31845e-39
	(b"10000000001100110101000011100100", b"00000000000000000000000000000000"),
	(b"00000000000110111101011100101010", b"10000000000101110111100110111010"), -- -4.71263e-39 + 2.55674e-39 = -2.15588e-39
	(b"00000000011100010011000101001111", b"00000000000000000000000000000000"),
	(b"00000000010110011001010011000000", b"00000000110010101100011000001111"), -- 1.03951e-38 + 8.22672e-39 = 1.86218e-38
	(b"00000000010000001001011000011111", b"00000000000000000000000000000000"),
	(b"00000000010000110010001110011010", b"00000000100000111011100110111001"), -- 5.93133e-39 + 6.16575e-39 = 1.20971e-38
	(b"10000000011011001110011011001011", b"00000000000000000000000000000000"),
	(b"00000000011001100001010111100100", b"10000000000001101101000011100111"), -- -1.0001e-38 + 9.37507e-39 = -6.25953e-40
	(b"10000000011011001110101111001001", b"00000000000000000000000000000000"),
	(b"10000000001001101100110000001010", b"10000000100100111011011111010011"), -- -1.00028e-38 + -3.56294e-39 = -1.35658e-38
	(b"00000000000111011101101011101100", b"00000000000000000000000000000000"),
	(b"00000000000000001111110111100000", b"00000000000111101101100011001100"), -- 2.74176e-39 + 9.10732e-41 = 2.83284e-39
	(b"10000000011000110000011000000111", b"00000000000000000000000000000000"),
	(b"00000000010110000110101111001001", b"10000000000010101001101000111110"), -- -9.09388e-39 + 8.12019e-39 = -9.73687e-40
	(b"10000000000011111100110000100001", b"00000000000000000000000000000000"),
	(b"00000000000000111110101011101001", b"10000000000010111110000100111000"), -- -1.45076e-39 + 3.59776e-40 = -1.09098e-39
	(b"10000000000100110111100010001011", b"00000000000000000000000000000000"),
	(b"00000000000100111101110011001100", b"00000000000000000110010001000001"), -- -1.78812e-39 + 1.82408e-39 = 3.59643e-41
	(b"10000000011001011110001101000000", b"00000000000000000000000000000000"),
	(b"10000000001001101000111001010000", b"10000000100011000111000110010000"), -- -9.35691e-39 + -3.5408e-39 = -1.28977e-38
	(b"00000000010101000110101110111100", b"00000000000000000000000000000000"),
	(b"00000000000010001101010110001010", b"00000000010111010100000101000110"), -- 7.75283e-39 + 8.11287e-40 = 8.56412e-39
	(b"10000000001011110011001110100010", b"00000000000000000000000000000000"),
	(b"10000000000100100000000010110111", b"10000000010000010011010001011001"), -- -4.33479e-39 + -1.6533e-39 = -5.98809e-39
	(b"10000000011011001101100100100111", b"00000000000000000000000000000000"),
	(b"10000000001010011010000001001001", b"10000000100101100111100101110000"), -- -9.99613e-39 + -3.82275e-39 = -1.38189e-38
	(b"00000000000010100111010111010110", b"00000000000000000000000000000000"),
	(b"00000000011110001010010001100111", b"00000000100000110001101000111101"), -- 9.60627e-40 + 1.10792e-38 = 1.20399e-38
	(b"10000000000010000010011100101111", b"00000000000000000000000000000000"),
	(b"00000000000000100100111111110011", b"10000000000001011101011100111100"), -- -7.4874e-40 + 2.12351e-40 = -5.36389e-40
	(b"00000000001111101000011011010000", b"00000000000000000000000000000000"),
	(b"00000000011110001010100000011010", b"00000000101101110010111011101010"), -- 5.74216e-39 + 1.10806e-38 = 1.68227e-38
	(b"00000000001111010011101010110000", b"00000000000000000000000000000000"),
	(b"00000000010100111011100000110011", b"00000000100100001111001011100011"), -- 5.62302e-39 + 7.68842e-39 = 1.33114e-38
	(b"00000000001000100101111011010110", b"00000000000000000000000000000000"),
	(b"10000000010011001000101111001010", b"10000000001010100010110011110100"), -- 3.15643e-39 + -7.02964e-39 = -3.87322e-39
	(b"10000000010011010101100101101111", b"00000000000000000000000000000000"),
	(b"00000000010011111011010010011011", b"00000000000000100101101100101100"), -- -7.10342e-39 + 7.31979e-39 = 2.16377e-40
	(b"00000000000011100010111000010101", b"00000000000000000000000000000000"),
	(b"00000000001010111010110011001101", b"00000000001110011101101011100010"), -- 1.30223e-39 + 4.01092e-39 = 5.31314e-39
	(b"10000000011100100100110101011011", b"00000000000000000000000000000000"),
	(b"00000000011100011111000100000010", b"10000000000000000101110001011001"), -- -1.0497e-38 + 1.04639e-38 = -3.31281e-41
	(b"10000000000101001110000001100100", b"00000000000000000000000000000000"),
	(b"00000000000010110110101100101011", b"10000000000010010111010100111001"), -- -1.91721e-39 + 1.04864e-39 = -8.68571e-40
	(b"10000000000111001010001011011011", b"00000000000000000000000000000000"),
	(b"00000000001110001101000101011001", b"00000000000111000010111001111110"), -- -2.62982e-39 + 5.21789e-39 = 2.58807e-39
	(b"00000000011000101010110010100011", b"00000000000000000000000000000000"),
	(b"00000000000010101101011010010001", b"00000000011011011000001100110100"), -- 9.06181e-39 + 9.95327e-40 = 1.00571e-38
	(b"10000000011110000101011001000000", b"00000000000000000000000000000000"),
	(b"10000000001001101000001111111110", b"10000000100111101101101000111110"), -- -1.10512e-38 + -3.5371e-39 = -1.45883e-38
	(b"00000000010010001100010100000101", b"00000000000000000000000000000000"),
	(b"10000000011000100110101000000011", b"10000000000110011010010011111110"), -- 6.68283e-39 + -9.03791e-39 = -2.35508e-39
	(b"10000000000011011010101000111010", b"00000000000000000000000000000000"),
	(b"00000000010001110110101101000111", b"00000000001110011100000100001101"), -- -1.25493e-39 + 6.5588e-39 = 5.30388e-39
	(b"00000000010110111011011011101011", b"00000000000000000000000000000000"),
	(b"00000000001010010101111100110110", b"00000000100001010001011000100001"), -- 8.42265e-39 + 3.79941e-39 = 1.22221e-38
	(b"10000000000000101111010100011000", b"00000000000000000000000000000000"),
	(b"10000000001001000111000011010010", b"10000000001001110110010111101010"), -- -2.71594e-40 + -3.34655e-39 = -3.61814e-39
	(b"00000000000011100110101111000101", b"00000000000000000000000000000000"),
	(b"00000000011111111010101101000100", b"00000000100011100001011100001001"), -- 1.32436e-39 + 1.17245e-38 = 1.30489e-38
	(b"10000000000100101010000010001010", b"00000000000000000000000000000000"),
	(b"10000000011100100010010101001001", b"10000000100001001100010111010011"), -- -1.71063e-39 + -1.04826e-38 = -1.21933e-38
	(b"00000000000110111001000011010110", b"00000000000000000000000000000000"),
	(b"00000000011001100110001010000010", b"00000000100000011111001101011000"), -- 2.53152e-39 + 9.40256e-39 = 1.19341e-38
	(b"10000000010100111110011111011011", b"00000000000000000000000000000000"),
	(b"10000000001001110010111100100000", b"10000000011110110001011011111011"), -- -7.70552e-39 + -3.59849e-39 = -1.1304e-38
	(b"10000000010111101100011101100000", b"00000000000000000000000000000000"),
	(b"00000000000000010100010110111111", b"10000000010111011000000110100001"), -- -8.70406e-39 + 1.16856e-40 = -8.5872e-39
	(b"00000000011101100011011111101110", b"00000000000000000000000000000000"),
	(b"00000000010110001101011001010110", b"00000000110011110000111001000100"), -- 1.08567e-38 + 8.15841e-39 = 1.90151e-38
	(b"10000000001111100010111011100110", b"00000000000000000000000000000000"),
	(b"10000000010101010100000010100010", b"10000000100100110110111110001000"), -- -5.71062e-39 + -7.8292e-39 = -1.35398e-38
	(b"00000000001010010100000001011000", b"00000000000000000000000000000000"),
	(b"00000000011111010010011111010001", b"00000000101001100110100000101001"), -- 3.78834e-39 + 1.14937e-38 = 1.52821e-38
	(b"00000000000101010101010110100110", b"00000000000000000000000000000000"),
	(b"10000000010011101010011010011100", b"10000000001110010101000011110110"), -- 1.95927e-39 + -7.22294e-39 = -5.26367e-39
	(b"00000000000100110000101101100110", b"00000000000000000000000000000000"),
	(b"00000000001010001110101110110010", b"00000000001110111111011100011000"), -- 1.74896e-39 + 3.75797e-39 = 5.50693e-39
	(b"10000000000011011011110001001001", b"00000000000000000000000000000000"),
	(b"10000000010111110011111000010000", b"10000000011011001111101001011001"), -- -1.26141e-39 + -8.74664e-39 = -1.0008e-38
	(b"10000000001111111000000111111101", b"00000000000000000000000000000000"),
	(b"10000000011000000000011001000110", b"10000000100111111000100001000011"), -- -5.83227e-39 + -8.81846e-39 = -1.46507e-38
	(b"10000000000111001001001100010000", b"00000000000000000000000000000000"),
	(b"00000000010101110010110100100010", b"00000000001110101001101000010010"), -- -2.62415e-39 + 8.00588e-39 = 5.38173e-39
	(b"00000000011110001010100001011000", b"00000000000000000000000000000000"),
	(b"00000000001001111100110011001101", b"00000000101000000111010100100101"), -- 1.10806e-38 + 3.65505e-39 = 1.47357e-38
	(b"00000000010001100110000010111001", b"00000000000000000000000000000000"),
	(b"00000000001011110011110111100100", b"00000000011101011001111010011101"), -- 6.46318e-39 + 4.33847e-39 = 1.08017e-38
	(b"10000000011111110111001110100101", b"00000000000000000000000000000000"),
	(b"00000000010000001100101101101011", b"10000000001111101010100000111010"), -- -1.17046e-38 + 5.95044e-39 = -5.75415e-39
	(b"10000000010111100010101011101010", b"00000000000000000000000000000000"),
	(b"00000000001011001000100011100110", b"10000000001100011010001000000100"), -- -8.64793e-39 + 4.08987e-39 = -4.55806e-39
	(b"00000000011110010110101110111010", b"00000000000000000000000000000000"),
	(b"00000000010101001100001000111000", b"00000000110011100010110111110010"), -- 1.11507e-38 + 7.78385e-39 = 1.89346e-38
	(b"10000000011011010000101011000110", b"00000000000000000000000000000000"),
	(b"00000000010101000000001110000110", b"10000000000110010000011101000000"), -- -1.00139e-38 + 7.71545e-39 = -2.29849e-39
	(b"00000000001101011111011011101000", b"00000000000000000000000000000000"),
	(b"10000000011101111111100110111010", b"10000000010000100000001011010010"), -- 4.95585e-39 + -1.1018e-38 = -6.06215e-39
	(b"10000000001010100110000111101101", b"00000000000000000000000000000000"),
	(b"10000000011000100111011000111101", b"10000000100011001101100000101010"), -- -3.89222e-39 + -9.04229e-39 = -1.29345e-38
	(b"00000000010111000010101010110110", b"00000000000000000000000000000000"),
	(b"10000000011101111110011101011101", b"10000000000110111011110010100111"), -- 8.46419e-39 + -1.10114e-38 = -2.54723e-39
	(b"00000000011010100001110110100011", b"00000000000000000000000000000000"),
	(b"10000000000101111101001011001111", b"00000000010100100100101011010100"), -- 9.74519e-39 + -2.18784e-39 = 7.55735e-39
	(b"10000000000100110001110100110100", b"00000000000000000000000000000000"),
	(b"00000000000110011001110100100000", b"00000000000001100111111111101100"), -- -1.75535e-39 + 2.35225e-39 = 5.96903e-40
	(b"00000000001100110111010100110100", b"00000000000000000000000000000000"),
	(b"00000000001010100011110011001011", b"00000000010111011011000111111111"), -- 4.72565e-39 + 3.8789e-39 = 8.60455e-39
	(b"10000000011100100010110001000101", b"00000000000000000000000000000000"),
	(b"10000000011111010101010101101010", b"10000000111011111000000110101111"), -- -1.04851e-38 + -1.15101e-38 = -2.19952e-38
	(b"00000000001111011110011101100001", b"00000000000000000000000000000000"),
	(b"10000000010011100110011100000011", b"10000000000100000111111110100010"), -- 5.68497e-39 + -7.20012e-39 = -1.51515e-39
	(b"00000000001001010000110110011101", b"00000000000000000000000000000000"),
	(b"10000000000001001100110011110010", b"00000000001000000100000010101011"), -- 3.4028e-39 + -4.40863e-40 = 2.96193e-39
	(b"10000000001101001010000010010011", b"00000000000000000000000000000000"),
	(b"10000000011100010100001111110000", b"10000000101001011110010010000011"), -- -4.83305e-39 + -1.04018e-38 = -1.52348e-38
	(b"00000000011100010111100100111001", b"00000000000000000000000000000000"),
	(b"00000000001011111100100011100101", b"00000000101000010100001000011110"), -- 1.04209e-38 + 4.38834e-39 = 1.48092e-38
	(b"10000000011110001001001011110001", b"00000000000000000000000000000000"),
	(b"00000000001100100010011110001011", b"10000000010001100110101101100110"), -- -1.1073e-38 + 4.60596e-39 = -6.46701e-39
	(b"00000000011110011110000110111111", b"00000000000000000000000000000000"),
	(b"10000000001011111011001000111110", b"00000000010010100010111110000001"), -- 1.11931e-38 + -4.38021e-39 = 6.81287e-39
	(b"10000000001001000111010101111111", b"00000000000000000000000000000000"),
	(b"00000000000111111111000110111110", b"10000000000001001000001111000001"), -- -3.34823e-39 + 2.93362e-39 = -4.14606e-40
	(b"10000000001000111001110011100110", b"00000000000000000000000000000000"),
	(b"10000000010011111101100100111101", b"10000000011100110111011000100011"), -- -3.27053e-39 + -7.33293e-39 = -1.06035e-38
	(b"10000000010111110000000000000111", b"00000000000000000000000000000000"),
	(b"10000000011010110011011000110011", b"10000000110010100011011000111010"), -- -8.72438e-39 + -9.84584e-39 = -1.85702e-38
	(b"00000000011010110101110000100100", b"00000000000000000000000000000000"),
	(b"00000000010000000100111010110001", b"00000000101010111010101011010101"), -- 9.85945e-39 + 5.9057e-39 = 1.57652e-38
	(b"10000000000001110010011000111000", b"00000000000000000000000000000000"),
	(b"00000000001100111011101111011110", b"00000000001011001001010110100110"), -- -6.56559e-40 + 4.751e-39 = 4.09445e-39
	(b"10000000010011011001001000000111", b"00000000000000000000000000000000"),
	(b"10000000000011010010100010110110", b"10000000010110101011101010111101"), -- -7.12372e-39 + -1.20847e-39 = -8.33218e-39
	(b"00000000001101100010001011001100", b"00000000000000000000000000000000"),
	(b"10000000000111100000110000010110", b"00000000000110000001011010110110"), -- 4.9716e-39 + -2.7594e-39 = 2.2122e-39
	(b"00000000010000011010011100000101", b"00000000000000000000000000000000"),
	(b"10000000010111001010110111101010", b"10000000000110110000011011100101"), -- 6.02922e-39 + -8.51125e-39 = -2.48203e-39
	(b"10000000011001111000101101001010", b"00000000000000000000000000000000"),
	(b"10000000001001101101011100101011", b"10000000100011100110001001110101"), -- -9.50902e-39 + -3.56694e-39 = -1.3076e-38
	(b"00000000000000111010111111110010", b"00000000000000000000000000000000"),
	(b"00000000000110110000111000000111", b"00000000000111101011110111111001"), -- 3.38624e-40 + 2.48459e-39 = 2.82321e-39
	(b"00000000001100101011111000001101", b"00000000000000000000000000000000"),
	(b"00000000000101011100110100000011", b"00000000010010001000101100010000"), -- 4.65995e-39 + 2.00209e-39 = 6.66204e-39
	(b"00000000001100010000001100101111", b"00000000000000000000000000000000"),
	(b"00000000000001100001001000001011", b"00000000001101110001010100111010"), -- 4.50108e-39 + 5.57486e-40 = 5.05857e-39
	(b"00000000000001010000000110101000", b"00000000000000000000000000000000"),
	(b"10000000010000111110100111001001", b"10000000001111101110100000100001"), -- 4.59772e-40 + -6.23684e-39 = -5.77707e-39
	(b"00000000000011001111010100101001", b"00000000000000000000000000000000"),
	(b"00000000001011110111100100011011", b"00000000001111000110111001000100"), -- 1.18997e-39 + 4.35971e-39 = 5.54969e-39
	(b"10000000001000110110100001011110", b"00000000000000000000000000000000"),
	(b"00000000010110110001101100001001", b"00000000001101111011001010101011"), -- -3.25168e-39 + 8.36673e-39 = 5.11505e-39
	(b"00000000001110010001101001001001", b"00000000000000000000000000000000"),
	(b"10000000000010001001101000000000", b"00000000001100001000000001001001"), -- 5.24405e-39 + -7.89929e-40 = 4.45412e-39
	(b"10000000001111001011100101000110", b"00000000000000000000000000000000"),
	(b"10000000011111000011011101100010", b"10000000101110001111000010101000"), -- -5.57659e-39 + -1.14075e-38 = -1.69841e-38
	(b"10000000000100000001111110000001", b"00000000000000000000000000000000"),
	(b"00000000010111101001101010110101", b"00000000010011100111101100110100"), -- -1.48067e-39 + 8.68804e-39 = 7.20737e-39
	(b"00000000001001011011111110111110", b"00000000000000000000000000000000"),
	(b"00000000011100000011101010000111", b"00000000100101011111101001000101"), -- 3.4667e-39 + 1.03066e-38 = 1.37733e-38
	(b"00000000001110011100111100000010", b"00000000000000000000000000000000"),
	(b"10000000001000111010100000111111", b"00000000000101100010011011000011"), -- 5.30888e-39 + -3.2746e-39 = 2.03429e-39
	(b"00000000001001010011100101101010", b"00000000000000000000000000000000"),
	(b"00000000011110100010011001101101", b"00000000100111110101111111010111"), -- 3.41851e-39 + 1.12177e-38 = 1.46362e-38
	(b"10000000001011011110111100011000", b"00000000000000000000000000000000"),
	(b"10000000000011000110001011011100", b"10000000001110100101000111110100"), -- -4.21837e-39 + -1.13749e-39 = -5.35586e-39
	(b"10000000001010111111101011010000", b"00000000000000000000000000000000"),
	(b"00000000001110001000101101100010", b"00000000000011001001000010010010"), -- -4.0389e-39 + 5.19279e-39 = 1.15389e-39
	(b"00000000000101011111001111000110", b"00000000000000000000000000000000"),
	(b"00000000010000111010010010000101", b"00000000010110011001100001001011"), -- 2.01599e-39 + 6.212e-39 = 8.22799e-39
	(b"10000000011111010111101010110000", b"00000000000000000000000000000000"),
	(b"10000000011010010101001011111000", b"10000000111001101100110110101000"), -- -1.15234e-38 + -9.67249e-39 = -2.11959e-38
	(b"10000000011011000000011001100010", b"00000000000000000000000000000000"),
	(b"00000000001001011101101110110100", b"10000000010001100010101010101110"), -- -9.92052e-39 + 3.47673e-39 = -6.4438e-39
	(b"00000000001000110100111001111011", b"00000000000000000000000000000000"),
	(b"10000000001010110000100111000100", b"10000000000001111011101101001001"), -- 3.2424e-39 + -3.95243e-39 = -7.10034e-40
	(b"10000000010110010100111110001010", b"00000000000000000000000000000000"),
	(b"00000000010110010111111100111110", b"00000000000000000010111110110100"), -- -8.20189e-39 + 8.21901e-39 = 1.71127e-41
	(b"10000000010000010101011000101111", b"00000000000000000000000000000000"),
	(b"00000000001100001000100000100110", b"10000000000100001100111000001001"), -- -6.00022e-39 + 4.45694e-39 = -1.54328e-39
	(b"00000000010111111011001010110000", b"00000000000000000000000000000000"),
	(b"10000000001011101011000010100110", b"00000000001100010000001000001010"), -- 8.78847e-39 + -4.2878e-39 = 4.50067e-39
	(b"10000000000100011110111010111111", b"00000000000000000000000000000000"),
	(b"10000000000110011101011110011101", b"10000000001010111100011001011100"), -- -1.64685e-39 + -2.37323e-39 = -4.02008e-39
	(b"00000000001111110001001100101100", b"00000000000000000000000000000000"),
	(b"00000000001000100110000000100110", b"00000000011000010111001101010010"), -- 5.79251e-39 + 3.1569e-39 = 8.94941e-39
	(b"10000000000100111000011101011000", b"00000000000000000000000000000000"),
	(b"10000000001101101011101010001100", b"10000000010010100100000111100100"), -- -1.79343e-39 + -5.02604e-39 = -6.81946e-39
	(b"10000000010010000010101111001000", b"00000000000000000000000000000000"),
	(b"10000000010001001101111101011000", b"10000000100011010000101100100000"), -- -6.62786e-39 + -6.32493e-39 = -1.29528e-38
	(b"00000000001010001001110110110010", b"00000000000000000000000000000000"),
	(b"00000000000010011000110100001100", b"00000000001100100010101010111110"), -- 3.72999e-39 + 8.77118e-40 = 4.60711e-39
	(b"10000000000101100000101111111001", b"00000000000000000000000000000000"),
	(b"10000000000001000111000101010111", b"10000000000110100111110101010000"), -- -2.02468e-39 + -4.08001e-40 = -2.43268e-39
	(b"10000000010010110000110111100011", b"00000000000000000000000000000000"),
	(b"00000000001101011001111000110111", b"10000000000101010110111110101100"), -- -6.89264e-39 + 4.92404e-39 = -1.96861e-39
	(b"00000000010010000101001010011110", b"00000000000000000000000000000000"),
	(b"10000000010011001101000101101001", b"10000000000001000111111011001011"), -- 6.64179e-39 + -7.05462e-39 = -4.12827e-40
	(b"00000000001111111011111101110000", b"00000000000000000000000000000000"),
	(b"10000000001010011111011001011100", b"00000000000101011100100100010100"), -- 5.85431e-39 + -3.85363e-39 = 2.00068e-39
	(b"00000000000111001100010110011000", b"00000000000000000000000000000000"),
	(b"00000000010011110111101111001010", b"00000000011011000100000101100010"), -- 2.64228e-39 + 7.29941e-39 = 9.94169e-39
	(b"10000000000101101110110110000110", b"00000000000000000000000000000000"),
	(b"10000000011011011011010101110110", b"10000000100001001010001011111100"), -- -2.10559e-39 + -1.00752e-38 = -1.21808e-38
	(b"10000000010101101010101110000001", b"00000000000000000000000000000000"),
	(b"00000000000001001001001100100000", b"10000000010100100001100001100001"), -- -7.95938e-39 + 4.2012e-40 = -7.53926e-39
	(b"00000000000010101100110100110011", b"00000000000000000000000000000000"),
	(b"00000000011100000001110011110101", b"00000000011110101110101000101000"), -- 9.91967e-40 + 1.0296e-38 = 1.12879e-38
	(b"00000000001010010101000110010111", b"00000000000000000000000000000000"),
	(b"10000000001101111101011100111111", b"10000000000011101000010110101000"), -- 3.79452e-39 + -5.12817e-39 = -1.33364e-39
	(b"10000000010110011111111010011010", b"00000000000000000000000000000000"),
	(b"10000000001101100000101110110001", b"10000000100100000000101001001011"), -- -8.26469e-39 + -4.96331e-39 = -1.3228e-38
	(b"00000000010110110001010010100001", b"00000000000000000000000000000000"),
	(b"00000000000111101100011100011101", b"00000000011110011101101110111110"), -- 8.36443e-39 + 2.82649e-39 = 1.11909e-38
	(b"00000000001100111010101110000011", b"00000000000000000000000000000000"),
	(b"00000000010010100000001101101001", b"00000000011111011010111011101100"), -- 4.74514e-39 + 6.79705e-39 = 1.15422e-38
	(b"10000000001101101111111001111010", b"00000000000000000000000000000000"),
	(b"00000000001000111110001110000111", b"10000000000100110001101011110011"), -- -5.05041e-39 + 3.29586e-39 = -1.75454e-39
	(b"10000000011001100010011111000100", b"00000000000000000000000000000000"),
	(b"10000000011010001011100100011101", b"10000000110011101110000011100001"), -- -9.38149e-39 + -9.6173e-39 = -1.89988e-38
	(b"10000000000001001101111111000100", b"00000000000000000000000000000000"),
	(b"10000000011111111110000110110100", b"10000000100001001100000101111000"), -- -4.47614e-40 + -1.17441e-38 = -1.21917e-38
	(b"00000000001100011100101010101001", b"00000000000000000000000000000000"),
	(b"00000000000111001111010001001011", b"00000000010011101011111011110100"), -- 4.57264e-39 + 2.65903e-39 = 7.23167e-39
	(b"10000000010110100000000000100010", b"00000000000000000000000000000000"),
	(b"00000000001101100110110000101111", b"10000000001000111001001111110011"), -- -8.26524e-39 + 4.99793e-39 = -3.26732e-39
	(b"10000000010010001000000111001101", b"00000000000000000000000000000000"),
	(b"00000000001010111001110100110001", b"10000000000111001110010010011100"), -- -6.65872e-39 + 4.00532e-39 = -2.6534e-39
	(b"10000000000100000110100110001001", b"00000000000000000000000000000000"),
	(b"00000000000010100010011110010111", b"10000000000001100100000111110010"), -- -1.50723e-39 + 9.32557e-40 = -5.7467e-40
	(b"00000000010001100110101110101111", b"00000000000000000000000000000000"),
	(b"10000000000010101110000111000111", b"00000000001110111000100111101000"), -- 6.46711e-39 + -9.99349e-40 = 5.46777e-39
	(b"00000000011000010110001100011111", b"00000000000000000000000000000000"),
	(b"10000000010101111010111010101011", b"00000000000010011011010001110100"), -- 8.9436e-39 + -8.05235e-39 = 8.91254e-40
	(b"00000000011100111111100001100101", b"00000000000000000000000000000000"),
	(b"00000000000110011101110111110100", b"00000000100011011101011001011001"), -- 1.06502e-38 + 2.37551e-39 = 1.30257e-38
	(b"00000000010011001101011111111101", b"00000000000000000000000000000000"),
	(b"00000000000010011110101000101000", b"00000000010101101100001000100101"), -- 7.05698e-39 + 9.10519e-40 = 7.9675e-39
	(b"10000000001110011011010001000101", b"00000000000000000000000000000000"),
	(b"10000000010110011010100010000011", b"10000000100100110101110011001000"), -- -5.29929e-39 + -8.23381e-39 = -1.35331e-38
	(b"00000000000100010100110111000110", b"00000000000000000000000000000000"),
	(b"10000000000101011110001010010111", b"10000000000001001001010011010001"), -- 1.5891e-39 + -2.00983e-39 = -4.20727e-40
	(b"10000000001011011111101100000011", b"00000000000000000000000000000000"),
	(b"10000000010110101110010100101010", b"10000000100010001110000000101101"), -- -4.22264e-39 + -8.3474e-39 = -1.257e-38
	(b"10000000010111001110101100001011", b"00000000000000000000000000000000"),
	(b"10000000000101100000100100000111", b"10000000011100101111010000010010"), -- -8.53318e-39 + -2.02362e-39 = -1.05568e-38
	(b"00000000010010011011010100101011", b"00000000000000000000000000000000"),
	(b"00000000010011000001010011100010", b"00000000100101011100101000001101"), -- 6.76898e-39 + 6.98699e-39 = 1.3756e-38
	(b"00000000011000010010111110101101", b"00000000000000000000000000000000"),
	(b"10000000010111100100101000011000", b"00000000000000101110010110010101"), -- 8.92515e-39 + -8.65912e-39 = 2.6603e-40
	(b"00000000000111111111000110110111", b"00000000000000000000000000000000"),
	(b"10000000000100011100010000011000", b"00000000000011100010110110011111"), -- 2.93361e-39 + -1.63155e-39 = 1.30206e-39
	(b"00000000010011101111100101001010", b"00000000000000000000000000000000"),
	(b"10000000010100000001111110101101", b"10000000000000010010011001100011"), -- 7.2526e-39 + -7.3582e-39 = -1.05606e-40
	(b"10000000000110011010101110111000", b"00000000000000000000000000000000"),
	(b"00000000001101000011101110000000", b"00000000000110101000111111001000"), -- -2.35749e-39 + 4.79679e-39 = 2.4393e-39
	(b"00000000010100001110110000001010", b"00000000000000000000000000000000"),
	(b"00000000000011100100010010100100", b"00000000010111110011000010101110"), -- 7.43151e-39 + 1.31032e-39 = 8.74184e-39
	(b"00000000011011110011101111010101", b"00000000000000000000000000000000"),
	(b"00000000011110000101100101110110", b"00000000111001111001010101001011"), -- 1.02152e-38 + 1.10524e-38 = 2.12676e-38
	(b"00000000001001001000111101100101", b"00000000000000000000000000000000"),
	(b"00000000000100010110000011000110", b"00000000001101011111000000101011"), -- 3.35752e-39 + 1.59592e-39 = 4.95344e-39
	(b"00000000000001110111110110001100", b"00000000000000000000000000000000"),
	(b"00000000001000101100111000010110", b"00000000001010100100101110100010"), -- 6.87886e-40 + 3.19634e-39 = 3.88422e-39
	(b"10000000000111011011000011110010", b"00000000000000000000000000000000"),
	(b"10000000010111001010100110010100", b"10000000011110100101101010000110"), -- -2.72671e-39 + -8.5097e-39 = -1.12364e-38
	(b"00000000000001111100100000001111", b"00000000000000000000000000000000"),
	(b"10000000001100011001001110101110", b"10000000001010011100101110011111"), -- 7.14616e-40 + -4.55292e-39 = -3.8383e-39
	(b"10000000011111111111001000011111", b"00000000000000000000000000000000"),
	(b"00000000001100111100100010100111", b"10000000010011000010100101111000"), -- -1.175e-38 + 4.75559e-39 = -6.99437e-39
	(b"10000000011110101110110001110101", b"00000000000000000000000000000000"),
	(b"10000000000100001010000010101011", b"10000000100010111000110100100000"), -- -1.12888e-38 + -1.527e-39 = -1.28158e-38
	(b"10000000010111100101011110110000", b"00000000000000000000000000000000"),
	(b"00000000010011011101111010111011", b"10000000000100000111100011110101"), -- -8.66399e-39 + 7.15123e-39 = -1.51276e-39
	(b"00000000010111101001111010010111", b"00000000000000000000000000000000"),
	(b"10000000000110110010101001100001", b"00000000010000110111010000110110"), -- 8.68943e-39 + -2.49476e-39 = 6.19467e-39
	(b"10000000001010001011110011100110", b"00000000000000000000000000000000"),
	(b"10000000000001001011100111101001", b"10000000001011010111011011001111"), -- -3.74118e-39 + -4.34034e-40 = -4.17522e-39
	(b"10000000011111110011111010010001", b"00000000000000000000000000000000"),
	(b"10000000001100101111100110101000", b"10000000101100100011100000111001"), -- -1.16856e-38 + -4.68133e-39 = -1.63669e-38
	(b"00000000001001101010010010010100", b"00000000000000000000000000000000"),
	(b"00000000001111100001101011110101", b"00000000011001001011111110001001"), -- 3.54879e-39 + 5.70347e-39 = 9.25226e-39
	(b"10000000000010001100000000010010", b"00000000000000000000000000000000"),
	(b"00000000011000101111111111110110", b"00000000010110100011111111100100"), -- -8.03586e-40 + 9.0917e-39 = 8.28811e-39
	(b"00000000010001100010000111100110", b"00000000000000000000000000000000"),
	(b"00000000001101010011000011111100", b"00000000011110110101001011100010"), -- 6.44065e-39 + 4.88485e-39 = 1.13255e-38
	(b"10000000001111010001011000110111", b"00000000000000000000000000000000"),
	(b"10000000010001010110111010001100", b"10000000100000101000010011000011"), -- -5.60993e-39 + -6.37631e-39 = -1.19862e-38
	(b"10000000000111000100001101110001", b"00000000000000000000000000000000"),
	(b"00000000001001100100110101100110", b"00000000000010100000100111110101"), -- -2.59559e-39 + 3.51751e-39 = 9.21927e-40
	(b"10000000000111101111010000100100", b"00000000000000000000000000000000"),
	(b"00000000011010001000101001001100", b"00000000010010011001011000101000"), -- -2.84265e-39 + 9.6005e-39 = 6.75786e-39
	(b"10000000001101100111010101101110", b"00000000000000000000000000000000"),
	(b"10000000001000011011111011000000", b"10000000010110000011010000101110"), -- -5.00124e-39 + -3.099e-39 = -8.10024e-39
	(b"00000000011001011101001110010011", b"00000000000000000000000000000000"),
	(b"00000000000010100001101001001011", b"00000000011011111110110111011110"), -- 9.35128e-39 + 9.27787e-40 = 1.02791e-38
	(b"10000000011001100001111011100111", b"00000000000000000000000000000000"),
	(b"10000000010100000110100011110011", b"10000000101101101000011111011010"), -- -9.37831e-39 + -7.38449e-39 = -1.67628e-38
	(b"10000000001101111000111000100101", b"00000000000000000000000000000000"),
	(b"00000000011101011110101101100110", b"00000000001111100101110101000001"), -- -5.10194e-39 + 1.08292e-38 = 5.72725e-39
	(b"00000000010101001101110010010011", b"00000000000000000000000000000000"),
	(b"10000000000101010011111111010100", b"00000000001111111001110010111111"), -- 7.79331e-39 + -1.95144e-39 = 5.84187e-39
	(b"00000000000101111011000011010011", b"00000000000000000000000000000000"),
	(b"10000000011111110011011000110101", b"10000000011001111000010101100010"), -- 2.17565e-39 + -1.16826e-38 = -9.5069e-39
	(b"10000000001110001100110101100010", b"00000000000000000000000000000000"),
	(b"00000000010010110101111100111100", b"00000000000100101001000111011010"), -- -5.21647e-39 + 6.92183e-39 = 1.70536e-39
	(b"00000000000010111111001100111110", b"00000000000000000000000000000000"),
	(b"10000000000011100000011101001000", b"10000000000000100001010000001010"), -- 1.09745e-39 + -1.28831e-39 = -1.9086e-40
	(b"00000000011100100000000111000110", b"00000000000000000000000000000000"),
	(b"00000000010100010100100011101001", b"00000000110000110100101010101111"), -- 1.04699e-38 + 7.46483e-39 = 1.79347e-38
	(b"00000000000011010111011111000011", b"00000000000000000000000000000000"),
	(b"00000000010010001100101111110101", b"00000000010101100100001110111000"), -- 1.23682e-39 + 6.68532e-39 = 7.92215e-39
	(b"10000000011011111011010101111101", b"00000000000000000000000000000000"),
	(b"10000000011100101110101010111111", b"10000000111000101010000000111100"), -- -1.02588e-38 + -1.05535e-38 = -2.08123e-38
	(b"10000000001110100010100110101100", b"00000000000000000000000000000000"),
	(b"10000000001111000100111001011000", b"10000000011101100111100000000100"), -- -5.34141e-39 + -5.53823e-39 = -1.08796e-38
	(b"00000000010001011001000100101011", b"00000000000000000000000000000000"),
	(b"10000000010010010100110000100100", b"10000000000000111011101011111001"), -- 6.38873e-39 + -6.73131e-39 = -3.4258e-40
	(b"10000000001100101001100001111101", b"00000000000000000000000000000000"),
	(b"10000000001001011100111010000011", b"10000000010110000110011100000000"), -- -4.64648e-39 + -3.472e-39 = -8.11847e-39
	(b"00000000010110101100001010001110", b"00000000000000000000000000000000"),
	(b"00000000011100001001010000010100", b"00000000110010110101011010100010"), -- 8.33499e-39 + 1.03387e-38 = 1.86737e-38
	(b"00000000011001000100000011100010", b"00000000000000000000000000000000"),
	(b"10000000011010100111101110011000", b"10000000000001100011101010110110"), -- 9.20683e-39 + -9.7789e-39 = -5.72074e-40
	(b"10000000001000110011101010010011", b"00000000000000000000000000000000"),
	(b"10000000000011001111101110000111", b"10000000001100000011011000011010"), -- -3.23525e-39 + -1.19226e-39 = -4.42751e-39
	(b"10000000000100001111000001100000", b"00000000000000000000000000000000"),
	(b"00000000000100011111011110101000", b"00000000000000010000011101001000"), -- -1.5556e-39 + 1.65005e-39 = 9.44475e-41
	(b"10000000011011001001000111110000", b"00000000000000000000000000000000"),
	(b"10000000000001001100010101000011", b"10000000011100010101011100110011"), -- -9.97059e-39 + -4.38106e-40 = -1.04087e-38
	(b"00000000011100000000110100110110", b"00000000000000000000000000000000"),
	(b"00000000010111111000011011101011", b"00000000110011111001010000100001"), -- 1.02903e-38 + 8.77277e-39 = 1.90631e-38
	(b"00000000010000010000111100011000", b"00000000000000000000000000000000"),
	(b"10000000000100101101101110101011", b"00000000001011100011001101101101"), -- 5.97472e-39 + -1.73184e-39 = 4.24288e-39
	(b"00000000000010110100011000010100", b"00000000000000000000000000000000"),
	(b"10000000011010100010101000011011", b"10000000010111101110010000000111"), -- 1.03533e-39 + -9.74967e-39 = -8.71434e-39
	(b"10000000000000111100101011101101", b"00000000000000000000000000000000"),
	(b"00000000010101110100011100101100", b"00000000010100110111110000111111"), -- -3.48303e-40 + 8.01522e-39 = 7.66692e-39
	(b"10000000011001010110000001011111", b"00000000000000000000000000000000"),
	(b"10000000000110110100100011100111", b"10000000100000001010100101000110"), -- -9.30996e-39 + -2.50571e-39 = -1.18157e-38
	(b"00000000001011010001011011111110", b"00000000000000000000000000000000"),
	(b"10000000010111000100100100000101", b"10000000001011110011001000000111"), -- 4.14085e-39 + -8.47506e-39 = -4.33421e-39
	(b"10000000001000000110100100000011", b"00000000000000000000000000000000"),
	(b"10000000001101011110101000111001", b"10000000010101100101001100111100"), -- -2.97641e-39 + -4.9513e-39 = -7.92771e-39
	(b"10000000011111101111101101101101", b"00000000000000000000000000000000"),
	(b"10000000010010001001100011001101", b"10000000110001111001010000111010"), -- -1.16615e-38 + -6.66697e-39 = -1.83284e-38
	(b"10000000001001011001101011101000", b"00000000000000000000000000000000"),
	(b"10000000011011100001011011000111", b"10000000100100111011000110101111"), -- -3.45348e-39 + -1.01101e-38 = -1.35636e-38
	(b"00000000001000111100010110110100", b"00000000000000000000000000000000"),
	(b"10000000000111010000111000101110", b"00000000000001101011011110000110"), -- 3.28516e-39 + -2.66832e-39 = 6.16849e-40
	(b"10000000010011001001111011000111", b"00000000000000000000000000000000"),
	(b"10000000000011000101110011101111", b"10000000010110001111101110110110"), -- -7.03646e-39 + -1.13536e-39 = -8.17182e-39
	(b"10000000010110010101111101011001", b"00000000000000000000000000000000"),
	(b"00000000000110000011011000110100", b"10000000010000010010100100100101"), -- -8.20756e-39 + 2.2235e-39 = -5.98407e-39
	(b"10000000000000000100110000100010", b"00000000000000000000000000000000"),
	(b"00000000010001101010011010010000", b"00000000010001100101101001101110"), -- -2.73113e-41 + 6.48824e-39 = 6.46092e-39
	(b"00000000001011001011001101111110", b"00000000000000000000000000000000"),
	(b"10000000011000011100001010010110", b"10000000001101010000111100011000"), -- 4.10515e-39 + -8.97785e-39 = -4.8727e-39
	(b"10000000000010001001011001110110", b"00000000000000000000000000000000"),
	(b"00000000000101000100101100110001", b"00000000000010111011010010111011"), -- -7.88659e-40 + 1.86368e-39 = 1.07502e-39
	(b"10000000011111110010101011100001", b"00000000000000000000000000000000"),
	(b"10000000000111110000101111000001", b"10000000100111100011011010100010"), -- -1.16785e-38 + -2.85112e-39 = -1.45296e-38
	(b"10000000000100011111010101011110", b"00000000000000000000000000000000"),
	(b"10000000001011001110100111001111", b"10000000001111101101111100101101"), -- -1.64922e-39 + -4.12464e-39 = -5.77386e-39
	(b"00000000000001001100011111110110", b"00000000000000000000000000000000"),
	(b"10000000000101101101011110100110", b"10000000000100100000111110110000"), -- 4.39074e-40 + -2.09774e-39 = -1.65867e-39
	(b"10000000011011000101001001111101", b"00000000000000000000000000000000"),
	(b"00000000010001000111000010011011", b"10000000001001111110000111100010"), -- -9.94782e-39 + 6.28521e-39 = -3.66262e-39
	(b"10000000000000001101011100001101", b"00000000000000000000000000000000"),
	(b"10000000001100011111110010011100", b"10000000001100101101001110101001"), -- -7.71457e-41 + -4.59056e-39 = -4.6677e-39
	(b"10000000010001000010010011101011", b"00000000000000000000000000000000"),
	(b"10000000001100101101101110010011", b"10000000011101110000000001111110"), -- -6.25806e-39 + -4.67054e-39 = -1.09286e-38
	(b"00000000000011111101001011011001", b"00000000000000000000000000000000"),
	(b"10000000011001000011010100000111", b"10000000010101000110001000101110"), -- 1.45317e-39 + -9.20257e-39 = -7.7494e-39
	(b"10000000010110000001110101100101", b"00000000000000000000000000000000"),
	(b"00000000011001100110011001001101", b"00000000000011100100100011101000"), -- -8.09207e-39 + 9.40392e-39 = 1.31185e-39
	(b"10000000000011100110001001011001", b"00000000000000000000000000000000"),
	(b"00000000001011010001111110111001", b"00000000000111101011110101100000"), -- -1.32098e-39 + 4.14398e-39 = 2.823e-39
	(b"10000000001011111000110100000011", b"00000000000000000000000000000000"),
	(b"10000000000001010100000000111010", b"10000000001101001100110100111101"), -- -4.36685e-39 + -4.82218e-40 = -4.84907e-39
	(b"00000000011110101001011101011010", b"00000000000000000000000000000000"),
	(b"00000000000100111110101000110010", b"00000000100011101000000110001100"), -- 1.12582e-38 + 1.82889e-39 = 1.30871e-38
	(b"10000000010001110101111001100100", b"00000000000000000000000000000000"),
	(b"00000000001000111000010010011001", b"10000000001000111101100111001011"), -- -6.55418e-39 + 3.26181e-39 = -3.29237e-39
	(b"10000000011000010110011111110000", b"00000000000000000000000000000000"),
	(b"00000000010110111111010011111000", b"10000000000001010111001011111000"), -- -8.94533e-39 + 8.44491e-39 = -5.0042e-40
	(b"00000000010010011101010000110100", b"00000000000000000000000000000000"),
	(b"10000000010010101110000101100010", b"10000000000000010000110100101110"), -- 6.78012e-39 + -6.87668e-39 = -9.65635e-41
	(b"10000000010010000011010110111001", b"00000000000000000000000000000000"),
	(b"00000000001000110001110101000100", b"10000000001001010001100001110101"), -- -6.63143e-39 + 3.22474e-39 = -3.40669e-39
	(b"00000000000011000000000100000101", b"00000000000000000000000000000000"),
	(b"10000000011110010101001111100010", b"10000000011011010101001011011101"), -- 1.10239e-39 + -1.11422e-38 = -1.00398e-38
	(b"00000000011111111001100111100100", b"00000000000000000000000000000000"),
	(b"00000000000011000110000000111110", b"00000000100010111111101000100010"), -- 1.17183e-38 + 1.13655e-39 = 1.28549e-38
	(b"10000000010110011000011111011110", b"00000000000000000000000000000000"),
	(b"10000000001010001011011010110011", b"10000000100000100011111010010001"), -- -8.2221e-39 + -3.73896e-39 = -1.19611e-38
	(b"10000000011010111100000010011010", b"00000000000000000000000000000000"),
	(b"00000000011001011011011001111100", b"10000000000001100000101000011110"), -- -9.89549e-39 + 9.34085e-39 = -5.54642e-40
	(b"00000000011000111110011110001111", b"00000000000000000000000000000000"),
	(b"00000000011001010000100010101101", b"00000000110010001111000000111100"), -- 9.17478e-39 + 9.2785e-39 = 1.84533e-38
	(b"10000000010010110000100101000111", b"00000000000000000000000000000000"),
	(b"00000000011001110000010110011100", b"00000000000110111111110001010101"), -- -6.89099e-39 + 9.46107e-39 = 2.57008e-39
	(b"00000000011111010100101000101101", b"00000000000000000000000000000000"),
	(b"00000000001000010010100010001010", b"00000000100111100111001010110111"), -- 1.1506e-38 + 3.04511e-39 = 1.45512e-38
	(b"10000000010111101111001111000011", b"00000000000000000000000000000000"),
	(b"10000000010000001011110101101110", b"10000000100111111011000100110001"), -- -8.71998e-39 + -5.94543e-39 = -1.46654e-38
	(b"00000000010001000001000110100100", b"00000000000000000000000000000000"),
	(b"00000000010110100110011110110100", b"00000000100111100111100101011000"), -- 6.25114e-39 + 8.3024e-39 = 1.45535e-38
	(b"10000000011110001100010100110000", b"00000000000000000000000000000000"),
	(b"00000000011101011011110111000011", b"10000000000000110000011101101101"), -- -1.1091e-38 + 1.08128e-38 = -2.7817e-40
	(b"00000000010100111111001010101101", b"00000000000000000000000000000000"),
	(b"00000000010101011111000011001000", b"00000000101010011110001101110101"), -- 7.7094e-39 + 7.89239e-39 = 1.56018e-38
	(b"00000000000011010100011001101000", b"00000000000000000000000000000000"),
	(b"10000000001011110100101001010001", b"10000000001000100000001111101001"), -- 1.21912e-39 + -4.34293e-39 = -3.12381e-39
	(b"10000000011101011011101001101111", b"00000000000000000000000000000000"),
	(b"00000000010011011000000100110000", b"10000000001010000011100100111111"), -- -1.08116e-38 + 7.11768e-39 = -3.69396e-39
	(b"00000000001010000011110010110111", b"00000000000000000000000000000000"),
	(b"10000000011100010000010100001001", b"10000000010010001100100001010010"), -- 3.6952e-39 + -1.03792e-38 = -6.68402e-39
	(b"00000000011000001001010100000001", b"00000000000000000000000000000000"),
	(b"10000000010101000101101110101000", b"00000000000011000011100101011001"), -- 8.86966e-39 + -7.74706e-39 = 1.1226e-39
	(b"10000000010011001111010010111101", b"00000000000000000000000000000000"),
	(b"10000000010100000000101010101100", b"10000000100111001111111101101001"), -- -7.06729e-39 + -7.35067e-39 = -1.4418e-38
	(b"10000000001001011110111101010001", b"00000000000000000000000000000000"),
	(b"10000000010101110111010011000001", b"10000000011111010110010000010010"), -- -3.48376e-39 + -8.03157e-39 = -1.15153e-38
	(b"00000000001010101000000111101000", b"00000000000000000000000000000000"),
	(b"10000000011100111101000111001000", b"10000000010010010100111111100000"), -- 3.90369e-39 + -1.06363e-38 = -6.73264e-39
	(b"10000000011000001000011010010100", b"00000000000000000000000000000000"),
	(b"10000000011010010000111010011000", b"10000000110010011001010100101100"), -- -8.86449e-39 + -9.64796e-39 = -1.85124e-38
	(b"10000000010010010100011011111010", b"00000000000000000000000000000000"),
	(b"00000000011110010100111100110000", b"00000000001100000000100000110110"), -- -6.72945e-39 + 1.11405e-38 = 4.41105e-39
	(b"00000000010000101010010101110000", b"00000000000000000000000000000000"),
	(b"10000000011111010001000111100101", b"10000000001110100110110001110101"), -- 6.12049e-39 + -1.14859e-38 = -5.36537e-39
	(b"00000000011110010111110000101111", b"00000000000000000000000000000000"),
	(b"10000000011011010111011100000000", b"00000000000011000000010100101111"), -- 1.11566e-38 + -1.00528e-38 = 1.10389e-39
	(b"00000000010100001100110100100000", b"00000000000000000000000000000000"),
	(b"10000000000111101010100011110111", b"00000000001100100010010000101001"), -- 7.42042e-39 + -2.81568e-39 = 4.60475e-39
	(b"10000000001111111101101011101110", b"00000000000000000000000000000000"),
	(b"10000000010011001110011101001010", b"10000000100011001100001000111000"), -- -5.86417e-39 + -7.06247e-39 = -1.29266e-38
	(b"00000000011011100000001010001101", b"00000000000000000000000000000000"),
	(b"10000000010011011100001000100100", b"00000000001000000100000001101001"), -- 1.01028e-38 + -7.14098e-39 = 2.96184e-39
	(b"00000000000110001010000010011010", b"00000000000000000000000000000000"),
	(b"10000000011110001100100000001010", b"10000000011000000010011101110000"), -- 2.26166e-39 + -1.1092e-38 = -8.83036e-39
	(b"10000000001101111011001101100010", b"00000000000000000000000000000000"),
	(b"00000000011000100000111100001110", b"00000000001010100101101110101100"), -- -5.1153e-39 + 9.00528e-39 = 3.88998e-39
	(b"10000000000010110110000000100001", b"00000000000000000000000000000000"),
	(b"10000000010100001111010111010011", b"10000000010111000101010111110100"), -- -1.04468e-39 + -7.43502e-39 = -8.4797e-39
	(b"00000000001101110011100111110111", b"00000000000000000000000000000000"),
	(b"00000000011011111100010011011011", b"00000000101001101111111011010010"), -- 5.07175e-39 + 1.02644e-38 = 1.53361e-38
	(b"00000000001001011101101010000101", b"00000000000000000000000000000000"),
	(b"00000000001100110011110000000000", b"00000000010110010001011010000101"), -- 3.4763e-39 + 4.70513e-39 = 8.18144e-39
	(b"10000000010010011010110010101111", b"00000000000000000000000000000000"),
	(b"10000000000110100000011100001000", b"10000000011000111011001110110111"), -- -6.76594e-39 + -2.39025e-39 = -9.15618e-39
	(b"10000000000110110111001111000111", b"00000000000000000000000000000000"),
	(b"00000000010101110001000111110001", b"00000000001110111001111000101010"), -- -2.52109e-39 + 7.99612e-39 = 5.47503e-39
	(b"00000000010000101111100100001110", b"00000000000000000000000000000000"),
	(b"10000000001110111000111100100110", b"00000000000001110110100111101000"), -- 6.15049e-39 + -5.46965e-39 = 6.8084e-40
	(b"10000000001000011011001110110001", b"00000000000000000000000000000000"),
	(b"00000000000010010101111000000100", b"10000000000110000101010110101101"), -- -3.09503e-39 + 8.60246e-40 = -2.23479e-39
	(b"10000000011110001010010110111001", b"00000000000000000000000000000000"),
	(b"00000000000110111110001010110010", b"10000000010111001100001100000111"), -- -1.10797e-38 + 2.56088e-39 = -8.51883e-39
	(b"00000000001111111010010011101101", b"00000000000000000000000000000000"),
	(b"10000000010001111111111111100011", b"10000000000010000101101011110110"), -- 5.8448e-39 + -6.61212e-39 = -7.67315e-40
	(b"00000000011010000100111100011101", b"00000000000000000000000000000000"),
	(b"00000000011010110001011010111111", b"00000000110100110110010111011100"), -- 9.57927e-39 + 9.83456e-39 = 1.94138e-38
	(b"00000000000011001101100011100111", b"00000000000000000000000000000000"),
	(b"10000000010101000111010001101110", b"10000000010001111001101110000111"), -- 1.17984e-39 + -7.75595e-39 = -6.57611e-39
	(b"00000000011111001010001110111110", b"00000000000000000000000000000000"),
	(b"10000000010101101011011010011110", b"00000000001001011110110100100000"), -- 1.14463e-38 + -7.96336e-39 = 3.48298e-39
	(b"10000000010010010011010000001001", b"00000000000000000000000000000000"),
	(b"00000000010000010100101011011111", b"10000000000001111110100100101010"), -- -6.72266e-39 + 5.99617e-39 = -7.26492e-40
	(b"00000000010110011100001001011000", b"00000000000000000000000000000000"),
	(b"10000000011100001110011010110101", b"10000000000101110010010001011101"), -- 8.24308e-39 + -1.03683e-38 = -2.12526e-39
	(b"10000000000001100000011000001010", b"00000000000000000000000000000000"),
	(b"10000000010111000010100101011001", b"10000000011000100010111101100011"), -- -5.53179e-40 + -8.4637e-39 = -9.01688e-39
	(b"00000000011001011010001101011111", b"00000000000000000000000000000000"),
	(b"10000000010000001100111100000111", b"00000000001001001101010001011000"), -- 9.33399e-39 + -5.95174e-39 = 3.38225e-39
	(b"00000000010000000001101011011110", b"00000000000000000000000000000000"),
	(b"00000000000010101110111100110000", b"00000000010010110000101000001110"), -- 5.88711e-39 + 1.00416e-39 = 6.89127e-39
	(b"00000000010100000010010000011000", b"00000000000000000000000000000000"),
	(b"00000000000100110010110111000010", b"00000000011000110101000111011010"), -- 7.35979e-39 + 1.76129e-39 = 9.12108e-39
	(b"10000000010110100100011110000010", b"00000000000000000000000000000000"),
	(b"00000000010100001011100011000011", b"10000000000010011000111010111111"), -- -8.29085e-39 + 7.41312e-39 = -8.77727e-40
	(b"00000000000110001110010011110100", b"00000000000000000000000000000000"),
	(b"10000000000011111001100101011101", b"00000000000010010100101110010111"), -- 2.28618e-39 + -1.43255e-39 = 8.53636e-40
	(b"10000000001010000110011011100000", b"00000000000000000000000000000000"),
	(b"00000000001001111001000101110110", b"10000000000000001101010101101010"), -- -3.71032e-39 + 3.63377e-39 = -7.65585e-41
	(b"10000000001111110001100001100100", b"00000000000000000000000000000000"),
	(b"00000000010101101011101010110001", b"00000000000101111010001001001101"), -- -5.79439e-39 + 7.96482e-39 = 2.17044e-39
	(b"00000000011000010000110100001001", b"00000000000000000000000000000000"),
	(b"10000000000010010101001010110000", b"00000000010101111011101001011001"), -- 8.91272e-39 + -8.56182e-40 = 8.05654e-39
	(b"00000000001111101010000010000001", b"00000000000000000000000000000000"),
	(b"10000000011100000101001100100011", b"10000000001100011011001010100010"), -- 5.75138e-39 + -1.03154e-38 = -4.56402e-39
	(b"00000000001000011001001100100001", b"00000000000000000000000000000000"),
	(b"10000000000010010110010110101010", b"00000000000110000010110101110111"), -- 3.08335e-39 + -8.6299e-40 = 2.22036e-39
	(b"00000000001011111110001010111001", b"00000000000000000000000000000000"),
	(b"00000000001110000100010010101010", b"00000000011010000010011101100011"), -- 4.3976e-39 + 5.16742e-39 = 9.56502e-39
	(b"00000000001111101101001010000110", b"00000000000000000000000000000000"),
	(b"00000000011111001011101010100101", b"00000000101110111000110100101011"), -- 5.76932e-39 + 1.14546e-38 = 1.72239e-38
	(b"00000000000011000000001000011101", b"00000000000000000000000000000000"),
	(b"00000000001010101101110001101000", b"00000000001101101101111010000101"), -- 1.10278e-39 + 3.93616e-39 = 5.03894e-39
	(b"10000000001001110010100111110101", b"00000000000000000000000000000000"),
	(b"00000000011110000011000110000010", b"00000000010100010000011110001101"), -- -3.59664e-39 + 1.1038e-38 = 7.44138e-39
	(b"00000000010111111001000110010010", b"00000000000000000000000000000000"),
	(b"10000000000011110100110101010101", b"00000000010100000100010000111101"), -- 8.77659e-39 + -1.40527e-39 = 7.37132e-39
	(b"00000000000001101010010010000100", b"00000000000000000000000000000000"),
	(b"00000000010000010010000111011001", b"00000000010001111100011001011101"), -- 6.1003e-40 + 5.98145e-39 = 6.59148e-39
	(b"10000000010101001001000100001001", b"00000000000000000000000000000000"),
	(b"10000000011101001010010010111000", b"10000000110010010011010111000001"), -- -7.76621e-39 + -1.0712e-38 = -1.84782e-38
	(b"10000000001001100101011011010000", b"00000000000000000000000000000000"),
	(b"00000000001110000101000100011100", b"00000000000100011111101001001100"), -- -3.52089e-39 + 5.17188e-39 = 1.65099e-39
	(b"00000000001101000001011011111101", b"00000000000000000000000000000000"),
	(b"00000000000110011001001011010101", b"00000000010011011010100111010010"), -- 4.78369e-39 + 2.34856e-39 = 7.13225e-39
	(b"00000000000001010100000011110111", b"00000000000000000000000000000000"),
	(b"10000000010111010100011011111110", b"10000000010110000000011000000111"), -- 4.82482e-40 + -8.56617e-39 = -8.08369e-39
	(b"00000000010011101001111110100001", b"00000000000000000000000000000000"),
	(b"00000000010010011001110110000111", b"00000000100110000011110100101000"), -- 7.22043e-39 + 6.7605e-39 = 1.39809e-38
	(b"00000000000000110110110111111100", b"00000000000000000000000000000000"),
	(b"00000000010000111100000000010111", b"00000000010001110010111000010011"), -- 3.14961e-40 + 6.22189e-39 = 6.53685e-39
	(b"10000000010100000010100001001010", b"00000000000000000000000000000000"),
	(b"10000000001110010011111000101001", b"10000000100010010110011001110011"), -- -7.36129e-39 + -5.25692e-39 = -1.26182e-38
	(b"10000000010010010000000000111000", b"00000000000000000000000000000000"),
	(b"00000000010111000100011101000110", b"00000000000100110100011100001110"), -- -6.70407e-39 + 8.47443e-39 = 1.77036e-39
	(b"00000000001010011101101000010000", b"00000000000000000000000000000000"),
	(b"00000000011100001010010111011110", b"00000000100110100111111111101110"), -- 3.84348e-39 + 1.03451e-38 = 1.41886e-38
	(b"00000000000110110111110101010011", b"00000000000000000000000000000000"),
	(b"00000000000101111110010000101100", b"00000000001100110110000101111111"), -- 2.52452e-39 + 2.19407e-39 = 4.71859e-39
	(b"10000000000000010111101101010011", b"00000000000000000000000000000000"),
	(b"10000000010111101101000100001000", b"10000000011000000100110001011011"), -- -1.36076e-40 + -8.70752e-39 = -8.8436e-39
	(b"10000000011111011100111110000001", b"00000000000000000000000000000000"),
	(b"00000000011011001010010100010010", b"10000000000100010010101001101111"), -- -1.15539e-38 + 9.97745e-39 = -1.57643e-39
	(b"10000000000010101011000110001101", b"00000000000000000000000000000000"),
	(b"00000000011101010110101110010010", b"00000000011010101011101000000101"), -- -9.82048e-40 + 1.07833e-38 = 9.80129e-39
	(b"00000000000101001100101110001101", b"00000000000000000000000000000000"),
	(b"10000000001110010001011110010011", b"10000000001001000100110000000110"), -- 1.90973e-39 + -5.24308e-39 = -3.33335e-39
	(b"10000000010100101111000100001111", b"00000000000000000000000000000000"),
	(b"10000000010011011111101000111110", b"10000000101000001110101101001101"), -- -7.61699e-39 + -7.1611e-39 = -1.47781e-38
	(b"00000000001100111000011010011011", b"00000000000000000000000000000000"),
	(b"00000000000111011110011111100010", b"00000000010100010110111001111101"), -- 4.7319e-39 + 2.74641e-39 = 7.47831e-39
	(b"00000000001011111001111011110111", b"00000000000000000000000000000000"),
	(b"00000000011011001010011110110010", b"00000000100111000100011010101001"), -- 4.37329e-39 + 9.97839e-39 = 1.43517e-38
	(b"10000000011010000001111011111010", b"00000000000000000000000000000000"),
	(b"00000000000110000101110100111111", b"10000000010011111100000110111011"), -- -9.562e-39 + 2.2375e-39 = -7.3245e-39
	(b"00000000011011010111010001011110", b"00000000000000000000000000000000"),
	(b"10000000010100000000011011010110", b"00000000000111010110110110001000"), -- 1.00518e-38 + -7.34929e-39 = 2.70252e-39
	(b"00000000010101001110001000010010", b"00000000000000000000000000000000"),
	(b"10000000010110011111010101010110", b"10000000000001010001001101000100"), -- 7.79528e-39 + -8.26137e-39 = -4.66089e-40
	(b"00000000001001101100000111100110", b"00000000000000000000000000000000"),
	(b"10000000000100010000100010110011", b"00000000000101011011100100110011"), -- 3.55931e-39 + -1.56432e-39 = 1.99498e-39
	(b"00000000001100110110100000111000", b"00000000000000000000000000000000"),
	(b"10000000010011010010011010011000", b"10000000000110011011111001100000"), -- 4.721e-39 + -7.08518e-39 = -2.36418e-39
	(b"10000000001000100110100110001111", b"00000000000000000000000000000000"),
	(b"00000000000011110000011001111011", b"10000000000100110110001100010100"), -- -3.16027e-39 + 1.37986e-39 = -1.78042e-39
	(b"10000000001111111100000110100001", b"00000000000000000000000000000000"),
	(b"10000000001111000001110010101010", b"10000000011110111101111001001011"), -- -5.8551e-39 + -5.52041e-39 = -1.13755e-38
	(b"10000000001100000100011001000110", b"00000000000000000000000000000000"),
	(b"00000000000101111000111100011010", b"10000000000110001011011100101100"), -- -4.43331e-39 + 2.16355e-39 = -2.26976e-39
	(b"10000000011000101010011110011011", b"00000000000000000000000000000000"),
	(b"10000000000110011011100100110000", b"10000000011111000110000011001011"), -- -9.06e-39 + -2.36232e-39 = -1.14223e-38
	(b"10000000010111011110001111100011", b"00000000000000000000000000000000"),
	(b"00000000010100011111001001001001", b"10000000000010111111000110011010"), -- -8.62245e-39 + 7.52559e-39 = -1.09686e-39
	(b"00000000011000101010001110001111", b"00000000000000000000000000000000"),
	(b"00000000011010000110000111101011", b"00000000110010110000010101111010"), -- 9.05855e-39 + 9.58602e-39 = 1.86446e-38
	(b"00000000011011000111111111100001", b"00000000000000000000000000000000"),
	(b"00000000011011111101101001111110", b"00000000110111000101101001011111"), -- 9.96411e-39 + 1.02721e-38 = 2.02362e-38
	(b"10000000000000110000010100111011", b"00000000000000000000000000000000"),
	(b"00000000001001110111100101001001", b"00000000001001000111010000001110"), -- -2.77383e-40 + 3.62509e-39 = 3.34771e-39
	(b"00000000010011101100000110000000", b"00000000000000000000000000000000"),
	(b"10000000001101010010111011110000", b"00000000000110011001001010010000"), -- 7.23258e-39 + -4.88412e-39 = 2.34846e-39
	(b"10000000001000011001011011111010", b"00000000000000000000000000000000"),
	(b"00000000001011011100101010101001", b"00000000000011000011001110101111"), -- -3.08473e-39 + 4.2053e-39 = 1.12057e-39
	(b"10000000010100010110111101011100", b"00000000000000000000000000000000"),
	(b"00000000001100001010110000010111", b"10000000001000001100001101000101"), -- -7.47862e-39 + 4.46984e-39 = -3.00879e-39
	(b"00000000000111100011001011100011", b"00000000000000000000000000000000"),
	(b"00000000010001010011110011010110", b"00000000011000110110111110111001"), -- 2.77332e-39 + 6.35847e-39 = 9.13179e-39
	(b"10000000010111000000110001100001", b"00000000000000000000000000000000"),
	(b"00000000001110111001010011111111", b"10000000001000000111011101100010"), -- -8.45331e-39 + 5.47174e-39 = -2.98156e-39
	(b"10000000010000111111000011100001", b"00000000000000000000000000000000"),
	(b"10000000000110100010010100000001", b"10000000010111100001010111100010"), -- -6.23939e-39 + -2.401e-39 = -8.64039e-39
	(b"10000000010010001111111000001000", b"00000000000000000000000000000000"),
	(b"10000000011101100111001011000101", b"10000000101111110111000011001101"), -- -6.70328e-39 + -1.08778e-38 = -1.7581e-38
	(b"10000000001010011100011100011101", b"00000000000000000000000000000000"),
	(b"10000000000010111010000010010101", b"10000000001101010110011110110010"), -- -3.83668e-39 + -1.0678e-39 = -4.90448e-39
	(b"10000000000100000111111000101101", b"00000000000000000000000000000000"),
	(b"10000000001100000000001010101000", b"10000000010000001000000011010101"), -- -1.51463e-39 + -4.40906e-39 = -5.92369e-39
	(b"00000000001010111001000100100011", b"00000000000000000000000000000000"),
	(b"00000000001001000000011000110111", b"00000000010011111001011101011010"), -- 4.00099e-39 + 3.30831e-39 = 7.3093e-39
	(b"10000000011011111100110000101101", b"00000000000000000000000000000000"),
	(b"00000000001110111100101111001111", b"10000000001101000000000001011110"), -- -1.0267e-38 + 5.49141e-39 = -4.77558e-39
	(b"10000000010111101000010111100101", b"00000000000000000000000000000000"),
	(b"10000000010101101000110011110001", b"10000000101101010001001011010110"), -- -8.68057e-39 + -7.94841e-39 = -1.6629e-38
	(b"10000000001010111010010000100111", b"00000000000000000000000000000000"),
	(b"10000000001001010100001000000011", b"10000000010100001110011000101010"), -- -4.00781e-39 + -3.42159e-39 = -7.42941e-39
	(b"00000000010011011101101010101101", b"00000000000000000000000000000000"),
	(b"00000000010111011000011001011010", b"00000000101010110110000100000111"), -- 7.14978e-39 + 8.5889e-39 = 1.57387e-38
	(b"10000000000101111111010101111110", b"00000000000000000000000000000000"),
	(b"00000000000001100110001010101100", b"10000000000100011001001011010010"), -- -2.20028e-39 + 5.8641e-40 = -1.61387e-39
	(b"10000000001001111001100001110111", b"00000000000000000000000000000000"),
	(b"10000000000001101010111010010111", b"10000000001011100100011100001110"), -- -3.63628e-39 + -6.13644e-40 = -4.24992e-39
	(b"10000000011111010001110101000010", b"00000000000000000000000000000000"),
	(b"10000000011110011110100110111010", b"10000000111101110000011011111100"), -- -1.14899e-38 + -1.11959e-38 = -2.26859e-38
	(b"00000000001111110011000011001000", b"00000000000000000000000000000000"),
	(b"00000000000010111000011011100111", b"00000000010010101011011110101111"), -- 5.80314e-39 + 1.05858e-39 = 6.86172e-39
	(b"10000000000011101011111111111000", b"00000000000000000000000000000000"),
	(b"00000000001001101100000010110010", b"00000000000110000000000010111010"), -- -1.35456e-39 + 3.55887e-39 = 2.20431e-39
	(b"10000000011100010101101101010110", b"00000000000000000000000000000000"),
	(b"00000000010001111100011110010000", b"10000000001010011001001111000110"), -- -1.04102e-38 + 6.59191e-39 = -3.81827e-39
	(b"10000000011001110001000001110010", b"00000000000000000000000000000000"),
	(b"00000000000001111011010001011001", b"10000000010111110101110000011001"), -- -9.46496e-39 + 7.07545e-40 = -8.75741e-39
	(b"10000000010000100111111001010000", b"00000000000000000000000000000000"),
	(b"00000000011011000111110100010110", b"00000000001010011111111011000110"), -- -6.10646e-39 + 9.96311e-39 = 3.85665e-39
	(b"00000000000011010100011010011011", b"00000000000000000000000000000000"),
	(b"10000000000001101111011110011000", b"00000000000001100100111100000011"), -- 1.21919e-39 + -6.39833e-40 = 5.79357e-40
	(b"10000000001011010000111010100011", b"00000000000000000000000000000000"),
	(b"10000000010001001000010001100111", b"10000000011100011001001100001010"), -- -4.13785e-39 + -6.29231e-39 = -1.04302e-38
	(b"10000000001101101111001001010101", b"00000000000000000000000000000000"),
	(b"10000000010011100001001011011111", b"10000000100001010000010100110100"), -- -5.04605e-39 + -7.16994e-39 = -1.2216e-38
	(b"00000000010010001001111100011011", b"00000000000000000000000000000000"),
	(b"10000000010011011010101100101011", b"10000000000001010000110000010000"), -- 6.66923e-39 + -7.13274e-39 = -4.63505e-40
	(b"00000000011000110001000100101000", b"00000000000000000000000000000000"),
	(b"00000000011011111111010101010010", b"00000000110100110000011001111010"), -- 9.09787e-39 + 1.02817e-38 = 1.93796e-38
	(b"10000000000111010100010001011101", b"00000000000000000000000000000000"),
	(b"00000000010000011111111101100010", b"00000000001001001011101100000101"), -- -2.68775e-39 + 6.06092e-39 = 3.37317e-39
	(b"10000000001111000011010110011111", b"00000000000000000000000000000000"),
	(b"10000000010001110110011010000011", b"10000000100000111001110000100010"), -- -5.52937e-39 + -6.55709e-39 = -1.20865e-38
	(b"10000000000110001111011011100110", b"00000000000000000000000000000000"),
	(b"00000000010011111011101110111001", b"00000000001101101100010011010011"), -- -2.29262e-39 + 7.32235e-39 = 5.02972e-39
	(b"00000000011000001101100110000110", b"00000000000000000000000000000000"),
	(b"00000000010110000100101001100001", b"00000000101110010010001111100111"), -- 8.89424e-39 + 8.10821e-39 = 1.70024e-38
	(b"10000000001010101001011110001101", b"00000000000000000000000000000000"),
	(b"10000000011011001100001001110001", b"10000000100101110101100111111110"), -- -3.91146e-39 + -9.98799e-39 = -1.38994e-38
	(b"00000000001101001001101110010111", b"00000000000000000000000000000000"),
	(b"10000000000100101010011110010111", b"00000000001000011111010000000000"), -- 4.83126e-39 + -1.71316e-39 = 3.1181e-39
	(b"00000000010100001010100010111010", b"00000000000000000000000000000000"),
	(b"10000000000011110111010100010111", b"00000000010000010011001110100011"), -- 7.40737e-39 + -1.41954e-39 = 5.98783e-39
	(b"00000000010001111001001011000100", b"00000000000000000000000000000000"),
	(b"10000000001000100000100100111100", b"00000000001001011000100110001000"), -- 6.57297e-39 + -3.12572e-39 = 3.44725e-39
	(b"00000000011010000101110000010010", b"00000000000000000000000000000000"),
	(b"10000000001011100110010011011110", b"00000000001110011111011100110100"), -- 9.58392e-39 + -4.26062e-39 = 5.3233e-39
	(b"00000000011110110100011100100011", b"00000000000000000000000000000000"),
	(b"00000000011110111110110001110101", b"00000000111101110011001110011000"), -- 1.13213e-38 + 1.13806e-38 = 2.27019e-38
	(b"00000000000001100111101010001110", b"00000000000000000000000000000000"),
	(b"10000000010001011111000101111000", b"10000000001111110111011011101010"), -- 5.94977e-40 + -6.42327e-39 = -5.82829e-39
	(b"10000000000101000010010001001010", b"00000000000000000000000000000000"),
	(b"10000000001010011110111010001011", b"10000000001111100001001011010101"), -- -1.84973e-39 + -3.85083e-39 = -5.70056e-39
	(b"10000000000010010100000000000110", b"00000000000000000000000000000000"),
	(b"00000000000101000001010001111110", b"00000000000010101101010001111000"), -- -8.49487e-40 + 1.84406e-39 = 9.94574e-40
	(b"00000000011010010001100101011000", b"00000000000000000000000000000000"),
	(b"00000000000011111101000110111101", b"00000000011110001110101100010101"), -- 9.65182e-39 + 1.45277e-39 = 1.11046e-38
	(b"10000000010110011001001111100111", b"00000000000000000000000000000000"),
	(b"10000000011011000110010101010111", b"10000000110001011111100100111110"), -- -8.22642e-39 + -9.95459e-39 = -1.8181e-38
	(b"10000000001010011010110001011010", b"00000000000000000000000000000000"),
	(b"00000000001001000110101111010000", b"10000000000001010100000010001010"), -- -3.82708e-39 + 3.34475e-39 = -4.8233e-40
	(b"00000000001111000111001001100000", b"00000000000000000000000000000000"),
	(b"10000000001011010101110100111110", b"00000000000011110001010100100010"), -- 5.55116e-39 + -4.16605e-39 = 1.38511e-39
	(b"00000000011010010110010001101000", b"00000000000000000000000000000000"),
	(b"00000000000111000110010101011010", b"00000000100001011100100111000010"), -- 9.67875e-39 + 2.60775e-39 = 1.22865e-38
	(b"10000000011111100111111000011010", b"00000000000000000000000000000000"),
	(b"10000000011101000111001110001110", b"10000000111100101111000110101000"), -- -1.16165e-38 + -1.06944e-38 = -2.23109e-38
	(b"00000000010001111111111101011011", b"00000000000000000000000000000000"),
	(b"00000000000100101011111001111110", b"00000000010110101011110111011001"), -- 6.61192e-39 + 1.72137e-39 = 8.3333e-39
	(b"10000000011001111101110111011010", b"00000000000000000000000000000000"),
	(b"10000000011111011010101111011010", b"10000000111001011000100110110100"), -- -9.53864e-39 + -1.15411e-38 = -2.10797e-38
	(b"00000000001101000101110000010101", b"00000000000000000000000000000000"),
	(b"10000000000011011111000011011000", b"00000000001001100110101100111101"), -- 4.80848e-39 + -1.28026e-39 = 3.52822e-39
	(b"00000000001100000001101010010001", b"00000000000000000000000000000000"),
	(b"10000000001111100001110010010001", b"10000000000011100000001000000000"), -- 4.41763e-39 + -5.70405e-39 = -1.28641e-39
	(b"00000000010011000110100101010000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000101100100", b"00000000010011000110011111101100"), -- 7.01728e-39 + -4.98862e-43 = 7.01678e-39
	(b"00000000000101101011001110001111", b"00000000000000000000000000000000"),
	(b"10000000000110001101011101101100", b"10000000000000100010001111011101"), -- 2.08479e-39 + -2.28133e-39 = -1.96536e-40
	(b"10000000011110111111111001010111", b"00000000000000000000000000000000"),
	(b"10000000010000111110100010011011", b"10000000101111111110011011110010"), -- -1.1387e-38 + -6.23642e-39 = -1.76234e-38
	(b"00000000011001110010000001010010", b"00000000000000000000000000000000"),
	(b"00000000000111000011001001001001", b"00000000100000110101001010011011"), -- 9.47065e-39 + 2.58943e-39 = 1.20601e-38
	(b"00000000000010100010011111100101", b"00000000000000000000000000000000"),
	(b"10000000011011100101110111100010", b"10000000011001000011010111111101"), -- 9.32666e-40 + -1.01356e-38 = -9.20292e-39
	(b"10000000000001100110010111000010", b"00000000000000000000000000000000"),
	(b"10000000010101111111100000010011", b"10000000010111100101110111010101"), -- -5.87517e-40 + -8.07868e-39 = -8.6662e-39
	(b"10000000011111010010100011100010", b"00000000000000000000000000000000"),
	(b"10000000011010011000001011010100", b"10000000111001101010101110110110"), -- -1.14941e-38 + -9.68966e-39 = -2.11838e-38
	(b"00000000000000000001110011110111", b"00000000000000000000000000000000"),
	(b"00000000011010110000011011110000", b"00000000011010110010001111100111"), -- 1.03906e-41 + 9.82889e-39 = 9.83928e-39
	(b"10000000011001001110100101110000", b"00000000000000000000000000000000"),
	(b"10000000010100111111101011110010", b"10000000101110001110010001100010"), -- -9.26729e-39 + -7.71237e-39 = -1.69797e-38
	(b"10000000010110000101110010001110", b"00000000000000000000000000000000"),
	(b"10000000011011110001101000010010", b"10000000110001110111011010100000"), -- -8.11473e-39 + -1.02031e-38 = -1.83178e-38
	(b"10000000011000000111111111100111", b"00000000000000000000000000000000"),
	(b"10000000001001010111101001001010", b"10000000100001011111101000110001"), -- -8.86209e-39 + -3.44178e-39 = -1.23039e-38
	(b"10000000010100001001000111010011", b"00000000000000000000000000000000"),
	(b"10000000010111110110100000000110", b"10000000101011111111100111011001"), -- -7.39915e-39 + -8.76169e-39 = -1.61608e-38
	(b"00000000001010010010011001000001", b"00000000000000000000000000000000"),
	(b"00000000001010110100101100001110", b"00000000010101000111000101001111"), -- 3.77898e-39 + 3.97585e-39 = 7.75483e-39
	(b"00000000010011101000010000110111", b"00000000000000000000000000000000"),
	(b"00000000011110100101011010100011", b"00000000110010001101101011011010"), -- 7.2106e-39 + 1.1235e-38 = 1.84456e-38
	(b"10000000010100001001010101000010", b"00000000000000000000000000000000"),
	(b"10000000011101111010011110000010", b"10000000110010000011110011000100"), -- -7.40038e-39 + -1.09885e-38 = -1.83889e-38
	(b"00000000001010001010110100101101", b"00000000000000000000000000000000"),
	(b"10000000000000010011110011010101", b"00000000001001110111000001011000"), -- 3.73554e-39 + -1.13658e-40 = 3.62189e-39
	(b"00000000000010110100111110010001", b"00000000000000000000000000000000"),
	(b"10000000000000000110001100011100", b"00000000000010101110110001110101"), -- 1.03873e-39 + -3.55537e-41 = 1.00318e-39
	(b"10000000011010111000111001011100", b"00000000000000000000000000000000"),
	(b"10000000001001001110101001101001", b"10000000100100000111100011000101"), -- -9.87747e-39 + -3.39017e-39 = -1.32676e-38
	(b"10000000011110010101001000010000", b"00000000000000000000000000000000"),
	(b"10000000001101110011111000101011", b"10000000101100001001000000111011"), -- -1.11415e-38 + -5.07325e-39 = -1.62148e-38
	(b"00000000011010001011101110101111", b"00000000000000000000000000000000"),
	(b"00000000001000100101010000010100", b"00000000100010110000111111000011"), -- 9.61822e-39 + 3.15257e-39 = 1.27708e-38
	(b"00000000011010011100111101111010", b"00000000000000000000000000000000"),
	(b"00000000001000000100011010011011", b"00000000100010100001011000010101"), -- 9.71716e-39 + 2.96406e-39 = 1.26812e-38
	(b"00000000000100001101111101010010", b"00000000000000000000000000000000"),
	(b"00000000011001101001100101000000", b"00000000011101110111100010010010"), -- 1.54948e-39 + 9.4222e-39 = 1.09717e-38
	(b"00000000011000001100010101101000", b"00000000000000000000000000000000"),
	(b"10000000001111011110100010111101", b"00000000001000101101110010101011"), -- 8.88702e-39 + -5.68546e-39 = 3.20157e-39
	(b"10000000001001101010110110010011", b"00000000000000000000000000000000"),
	(b"10000000001111101101000000000101", b"10000000011001010111110110011000"), -- -3.55202e-39 + -5.76842e-39 = -9.32044e-39
	(b"10000000001011101111000001000111", b"00000000000000000000000000000000"),
	(b"10000000010011110100110001011000", b"10000000011111100011110010011111"), -- -4.31063e-39 + -7.28239e-39 = -1.1593e-38
	(b"00000000000000100110010000001001", b"00000000000000000000000000000000"),
	(b"00000000000010101110010101101000", b"00000000000011010100100101110001"), -- 2.19557e-40 + 1.00065e-39 = 1.22021e-39
	(b"10000000011100001010010101101011", b"00000000000000000000000000000000"),
	(b"00000000010011000101110110000111", b"10000000001001000100011111100100"), -- -1.03449e-38 + 7.01305e-39 = -3.33187e-39
	(b"00000000001101111111010010110010", b"00000000000000000000000000000000"),
	(b"00000000001000011001110100101110", b"00000000010110011001000111100000"), -- 5.13873e-39 + 3.08696e-39 = 8.22569e-39
	(b"10000000001111100111110010010100", b"00000000000000000000000000000000"),
	(b"00000000010111000110100110100111", b"00000000000111011110110100010011"), -- -5.73849e-39 + 8.48677e-39 = 2.74828e-39
	(b"00000000001111000001001001111111", b"00000000000000000000000000000000"),
	(b"10000000001001001010100110001101", b"00000000000101110110100011110010"), -- 5.51676e-39 + -3.3669e-39 = 2.14986e-39
	(b"00000000010100110010011100000101", b"00000000000000000000000000000000"),
	(b"10000000000000010100110110000110", b"00000000010100011101100101111111"), -- 7.63634e-39 + -1.19646e-40 = 7.5167e-39
	(b"10000000001111000111111111110100", b"00000000000000000000000000000000"),
	(b"00000000011110110101010111011000", b"00000000001111101101010111100100"), -- -5.55603e-39 + 1.13266e-38 = 5.77053e-39
	(b"00000000011101100110010011101011", b"00000000000000000000000000000000"),
	(b"00000000001111100010101110101101", b"00000000101101001001000010011000"), -- 1.08728e-38 + 5.70947e-39 = 1.65823e-38
	(b"00000000000100111011100110110101", b"00000000000000000000000000000000"),
	(b"00000000010100010110000010011101", b"00000000011001010001101001010010"), -- 1.81149e-39 + 7.47333e-39 = 9.28483e-39
	(b"10000000000111111001110001001011", b"00000000000000000000000000000000"),
	(b"00000000010110001101000111111000", b"00000000001110010011010110101101"), -- -2.90297e-39 + 8.15685e-39 = 5.25388e-39
	(b"10000000010011001000011000001011", b"00000000000000000000000000000000"),
	(b"10000000001011001100100000100101", b"10000000011110010100111000110000"), -- -7.02758e-39 + -4.11256e-39 = -1.11401e-38
	(b"00000000000111001101111000000100", b"00000000000000000000000000000000"),
	(b"00000000010100001010110111000010", b"00000000011011011000101111000110"), -- 2.65104e-39 + 7.40917e-39 = 1.00602e-38
	(b"00000000010110100010101110111010", b"00000000000000000000000000000000"),
	(b"00000000001101111110111100000000", b"00000000100100100001101010111010"), -- 8.28088e-39 + 5.13669e-39 = 1.34176e-38
	(b"00000000010100010111110010001001", b"00000000000000000000000000000000"),
	(b"10000000011011110000110100101010", b"10000000000111011001000010100001"), -- 7.48335e-39 + -1.01985e-38 = -2.71511e-39
	(b"10000000001111110100010110010100", b"00000000000000000000000000000000"),
	(b"00000000011001010001111011011011", b"00000000001001011101100101000111"), -- -5.8106e-39 + 9.28645e-39 = 3.47586e-39
	(b"10000000011110111100100100000111", b"00000000000000000000000000000000"),
	(b"10000000000100011100101110011110", b"10000000100011011001010010100101"), -- -1.13679e-38 + -1.63425e-39 = -1.30021e-38
	(b"10000000010000101010101000011111", b"00000000000000000000000000000000"),
	(b"00000000000000111101000001100100", b"10000000001111101101100110111011"), -- -6.12217e-39 + 3.50263e-40 = -5.77191e-39
	(b"10000000001101101011100010100101", b"00000000000000000000000000000000"),
	(b"00000000000000010111111110000111", b"10000000001101010011100100011110"), -- -5.02535e-39 + 1.37584e-40 = -4.88777e-39
	(b"00000000001100011101110100001000", b"00000000000000000000000000000000"),
	(b"00000000010111110001001100111000", b"00000000100100001111000001000000"), -- 4.57923e-39 + 8.73127e-39 = 1.33105e-38
	(b"10000000001101010011001111100011", b"00000000000000000000000000000000"),
	(b"10000000010110011110100100101101", b"10000000100011110001110100010000"), -- -4.88589e-39 + -8.25701e-39 = -1.31429e-38
	(b"00000000010010001100101011001111", b"00000000000000000000000000000000"),
	(b"00000000011000011111110101111111", b"00000000101010101100100001001110"), -- 6.68491e-39 + 8.99898e-39 = 1.56839e-38
	(b"10000000000111001111001001101000", b"00000000000000000000000000000000"),
	(b"00000000011000101100100110001111", b"00000000010001011101011100100111"), -- -2.65835e-39 + 9.07218e-39 = 6.41383e-39
	(b"00000000010110101010001111000001", b"00000000000000000000000000000000"),
	(b"00000000001000001010001101110011", b"00000000011110110100011100110100"), -- 8.32394e-39 + 2.99737e-39 = 1.13213e-38
	(b"10000000000101011110001000110001", b"00000000000000000000000000000000"),
	(b"10000000001110110100011101101010", b"10000000010100010010100110011011"), -- -2.00969e-39 + -5.44391e-39 = -7.4536e-39
	(b"10000000011000010001100111011011", b"00000000000000000000000000000000"),
	(b"00000000000001001011010010010100", b"10000000010111000110010101000111"), -- -8.91732e-39 + 4.32121e-40 = -8.4852e-39
	(b"00000000000101010011001101000001", b"00000000000000000000000000000000"),
	(b"10000000000011010110110101110101", b"00000000000001111100010111001100"), -- 1.94693e-39 + -1.23313e-39 = 7.13805e-40
	(b"00000000010011110010110011111111", b"00000000000000000000000000000000"),
	(b"00000000000100100011111011111000", b"00000000011000010110101111110111"), -- 7.27115e-39 + 1.67563e-39 = 8.94677e-39
	(b"00000000001111011000111011001111", b"00000000000000000000000000000000"),
	(b"10000000000000010100000111001011", b"00000000001111000100110100000100"), -- 5.6532e-39 + -1.15438e-40 = 5.53776e-39
	(b"10000000011111101101010110001101", b"00000000000000000000000000000000"),
	(b"00000000011001001001111010010111", b"10000000000110100011011011110110"), -- -1.16479e-38 + 9.24044e-39 = -2.40744e-39
	(b"10000000001001000110000011010111", b"00000000000000000000000000000000"),
	(b"10000000001111100001010100010101", b"10000000011000100111010111101100"), -- -3.34082e-39 + -5.70136e-39 = -9.04218e-39
	(b"10000000001001101101110011111011", b"00000000000000000000000000000000"),
	(b"00000000000001011110100000001111", b"10000000001000001111010011101100"), -- -3.56902e-39 + 5.42424e-40 = -3.0266e-39
	(b"00000000001101101111101000011011", b"00000000000000000000000000000000"),
	(b"10000000001110111100010110111100", b"10000000000001001100101110100001"), -- 5.04884e-39 + -5.48923e-39 = -4.4039e-40
	(b"00000000001000110010100110011100", b"00000000000000000000000000000000"),
	(b"00000000011100000000101110010001", b"00000000100100110011010100101101"), -- 3.22917e-39 + 1.02897e-38 = 1.35189e-38
	(b"00000000010010010110011101101101", b"00000000000000000000000000000000"),
	(b"00000000001100111100010111011010", b"00000000011111010010110101000111"), -- 6.74109e-39 + 4.75459e-39 = 1.14957e-38
	(b"00000000011000111110011100110111", b"00000000000000000000000000000000"),
	(b"00000000010000101001101010001000", b"00000000101001101000000110111111"), -- 9.17466e-39 + 6.11658e-39 = 1.52912e-38
	(b"10000000010111101010100110110110", b"00000000000000000000000000000000"),
	(b"00000000001101000010010110010000", b"10000000001010101000010000100110"), -- -8.69342e-39 + 4.78892e-39 = -3.9045e-39
	(b"00000000010101010110100010000111", b"00000000000000000000000000000000"),
	(b"10000000000110011111100111001011", b"00000000001110110110111010111100"), -- 7.84351e-39 + -2.3855e-39 = 5.45802e-39
	(b"00000000001011100001110100001000", b"00000000000000000000000000000000"),
	(b"00000000001111100011011011010110", b"00000000011011000101001111011110"), -- 4.23485e-39 + 5.71347e-39 = 9.94832e-39
	(b"10000000011000100010011011111100", b"00000000000000000000000000000000"),
	(b"10000000010011111100100110010111", b"10000000101100011111000010010011"), -- -9.01386e-39 + -7.32732e-39 = -1.63412e-38
	(b"10000000010101001111101110111100", b"00000000000000000000000000000000"),
	(b"10000000010010011111001011011010", b"10000000100111101110111010010110"), -- -7.80449e-39 + -6.79111e-39 = -1.45956e-38
	(b"00000000001001001011100100100000", b"00000000000000000000000000000000"),
	(b"00000000000011010001001101001111", b"00000000001100011100110001101111"), -- 3.37249e-39 + 1.20079e-39 = 4.57328e-39
	(b"00000000000011010011000011001010", b"00000000000000000000000000000000"),
	(b"00000000001111111111101100001001", b"00000000010011010010101111010011"), -- 1.21136e-39 + 5.87569e-39 = 7.08705e-39
	(b"00000000000010100110000101101001", b"00000000000000000000000000000000"),
	(b"10000000011110011111111001011000", b"10000000011011111001110011101111"), -- 9.53299e-40 + -1.12033e-38 = -1.025e-38
	(b"10000000000111110001011011110001", b"00000000000000000000000000000000"),
	(b"00000000010100101110001010110011", b"00000000001100111100101111000010"), -- -2.85513e-39 + 7.61184e-39 = 4.7567e-39
	(b"00000000011100000100010101011011", b"00000000000000000000000000000000"),
	(b"00000000000010001000101110010010", b"00000000011110001101000011101101"), -- 1.03105e-38 + 7.84752e-40 = 1.10952e-38
	(b"00000000001110111001111101010100", b"00000000000000000000000000000000"),
	(b"00000000001000000010010100111101", b"00000000010110111100010010010001"), -- 5.47545e-39 + 2.95209e-39 = 8.42754e-39
	(b"00000000000110101111001101101000", b"00000000000000000000000000000000"),
	(b"10000000000100011101110010010000", b"00000000000010010001011011011000"), -- 2.47504e-39 + -1.64033e-39 = 8.34714e-40
	(b"10000000011101101011010100100011", b"00000000000000000000000000000000"),
	(b"00000000000110000000100111000111", b"10000000010111101010101101011100"), -- -1.09016e-38 + 2.20756e-39 = -8.69401e-39
	(b"10000000011010000010110011101101", b"00000000000000000000000000000000"),
	(b"00000000001101101011011110011010", b"10000000001100010111010101010011"), -- -9.56701e-39 + 5.02498e-39 = -4.54203e-39
	(b"00000000001110001111110111000001", b"00000000000000000000000000000000"),
	(b"00000000010001100101001101010001", b"00000000011111110101000100010010"), -- 5.23382e-39 + 6.45837e-39 = 1.16922e-38
	(b"00000000000110101101011101101001", b"00000000000000000000000000000000"),
	(b"00000000010100110010110001000100", b"00000000011011100000001110101101"), -- 2.465e-39 + 7.63823e-39 = 1.01032e-38
	(b"00000000001011010100110010111101", b"00000000000000000000000000000000"),
	(b"00000000001001101001001101111101", b"00000000010100111110000000111010"), -- 4.16013e-39 + 3.54266e-39 = 7.70278e-39
	(b"10000000011100001111001100111010", b"00000000000000000000000000000000"),
	(b"00000000011101000011110001001010", b"00000000000000110100100100010000"), -- -1.03728e-38 + 1.06745e-38 = 3.01716e-40
	(b"10000000010100110111000000111111", b"00000000000000000000000000000000"),
	(b"00000000001011100001101001100110", b"10000000001001010101010111011001"), -- -7.66261e-39 + 4.2339e-39 = -3.42871e-39
	(b"10000000011011100100111000000100", b"00000000000000000000000000000000"),
	(b"10000000010110110010100010011011", b"10000000110010010111011010011111"), -- -1.01299e-38 + -8.3716e-39 = -1.85015e-38
	(b"00000000001001101011011010010000", b"00000000000000000000000000000000"),
	(b"00000000011010110100001000010010", b"00000000100100011111100010100010"), -- 3.55524e-39 + 9.8501e-39 = 1.34053e-38
	(b"10000000010101010010110100011000", b"00000000000000000000000000000000"),
	(b"10000000000111111101000110110100", b"10000000011101001111111011001100"), -- -7.82219e-39 + -2.92213e-39 = -1.07443e-38
	(b"00000000011111001100000110110101", b"00000000000000000000000000000000"),
	(b"10000000010001000011010101010111", b"00000000001110001000110001011110"), -- 1.14571e-38 + -6.26395e-39 = 5.19314e-39
	(b"10000000010101101101010011100110", b"00000000000000000000000000000000"),
	(b"10000000000101011011011010110010", b"10000000011011001000101110011000"), -- -7.97423e-39 + -1.99408e-39 = -9.96831e-39
	(b"10000000000101000111101011010111", b"00000000000000000000000000000000"),
	(b"10000000001010010001010011011000", b"10000000001111011000111110101111"), -- -1.88078e-39 + -3.77273e-39 = -5.65351e-39
	(b"00000000000011010011101000001110", b"00000000000000000000000000000000"),
	(b"00000000010101011000101000001110", b"00000000011000101100010000011100"), -- 1.21469e-39 + 7.85554e-39 = 9.07023e-39
	(b"10000000010011101001000010001101", b"00000000000000000000000000000000"),
	(b"00000000001000001101000011111100", b"10000000001011011011111110010001"), -- -7.21502e-39 + 3.01371e-39 = -4.20132e-39
	(b"00000000011100110111011010100001", b"00000000000000000000000000000000"),
	(b"00000000001110111010111110111100", b"00000000101011110010011001011101"), -- 1.06036e-38 + 5.48134e-39 = 1.6085e-38
	(b"10000000000100101001100010010000", b"00000000000000000000000000000000"),
	(b"10000000010000101011010001000100", b"10000000010101010100110011010100"), -- -1.70777e-39 + -6.12581e-39 = -7.83358e-39
	(b"00000000001101001101010011101110", b"00000000000000000000000000000000"),
	(b"00000000000000010010101010101100", b"00000000001101011111111110011010"), -- 4.85183e-39 + 1.07143e-40 = 4.95897e-39
	(b"00000000010100011101111011010001", b"00000000000000000000000000000000"),
	(b"00000000011011111011001011101010", b"00000000110000011001000110111011"), -- 7.51861e-39 + 1.02579e-38 = 1.77765e-38
	(b"10000000011100000001111101000111", b"00000000000000000000000000000000"),
	(b"10000000010011000001100001101100", b"10000000101111000011011110110011"), -- -1.02968e-38 + -6.98826e-39 = -1.72851e-38
	(b"10000000010101000101111101010110", b"00000000000000000000000000000000"),
	(b"00000000001000000100010110000110", b"10000000001101000001100111010000"), -- -7.74838e-39 + 2.96368e-39 = -4.78471e-39
	(b"10000000010100110011001111000010", b"00000000000000000000000000000000"),
	(b"10000000000111101001110111001010", b"10000000011100011101000110001100"), -- -7.64091e-39 + -2.81167e-39 = -1.04526e-38
	(b"00000000000100110100100010111111", b"00000000000000000000000000000000"),
	(b"10000000001111010111010100010101", b"10000000001010100010110001010110"), -- 1.77097e-39 + -5.64397e-39 = -3.873e-39
	(b"10000000011000110101100101000100", b"00000000000000000000000000000000"),
	(b"10000000010011010101110010000110", b"10000000101100001011010111001010"), -- -9.12374e-39 + -7.10452e-39 = -1.62283e-38
	(b"10000000010001101100011111111000", b"00000000000000000000000000000000"),
	(b"10000000010011010001010110101000", b"10000000100100111101110110100000"), -- -6.50022e-39 + -7.0791e-39 = -1.35793e-38
	(b"00000000001011011011110001111110", b"00000000000000000000000000000000"),
	(b"10000000001110100110000000010000", b"10000000000011001010001110010010"), -- 4.20022e-39 + -5.36092e-39 = -1.1607e-39
	(b"00000000000010111000000101001001", b"00000000000000000000000000000000"),
	(b"00000000011100000111101011000001", b"00000000011110111111110000001010"), -- 1.05657e-39 + 1.03296e-38 = 1.13862e-38
	(b"10000000000010100100010011111000", b"00000000000000000000000000000000"),
	(b"00000000010010000111111001000110", b"00000000001111100011100101001110"), -- -9.43096e-40 + 6.65745e-39 = 5.71436e-39
	(b"10000000000101100111111110111000", b"00000000000000000000000000000000"),
	(b"00000000000100110101011001111110", b"10000000000000110010100100111010"), -- -2.0662e-39 + 1.7759e-39 = -2.90296e-40
	(b"10000000011000001010111011000110", b"00000000000000000000000000000000"),
	(b"00000000000111110011110010010110", b"10000000010000010111001000110000"), -- -8.8789e-39 + 2.86863e-39 = -6.01027e-39
	(b"00000000011110101100101011010000", b"00000000000000000000000000000000"),
	(b"10000000000101001000000100011111", b"00000000011001100100100110110001"), -- 1.12767e-38 + -1.88303e-39 = 9.39366e-39
	(b"00000000000101101001001011111100", b"00000000000000000000000000000000"),
	(b"00000000011111111100011100010001", b"00000000100101100101101000001101"), -- 2.07311e-39 + 1.17345e-38 = 1.38076e-38
	(b"10000000011111101111111100001010", b"00000000000000000000000000000000"),
	(b"10000000000111001101010100001001", b"10000000100110111101010000010011"), -- -1.16628e-38 + -2.64782e-39 = -1.43106e-38
	(b"00000000001110010111001111101011", b"00000000000000000000000000000000"),
	(b"00000000011011010101000101001100", b"00000000101001101100010100110111"), -- 5.27621e-39 + 1.00392e-38 = 1.53154e-38
	(b"10000000010100111110101001110110", b"00000000000000000000000000000000"),
	(b"00000000000110101010110101001111", b"10000000001110010011110100100111"), -- -7.70645e-39 + 2.44989e-39 = -5.25656e-39
	(b"00000000000000000011101010101110", b"00000000000000000000000000000000"),
	(b"00000000011001111010010011100111", b"00000000011001111101111110010101"), -- 2.10503e-41 + 9.51821e-39 = 9.53926e-39
	(b"00000000001000000011100100101000", b"00000000000000000000000000000000"),
	(b"10000000010010000011110110001111", b"10000000001010000000010001100111"), -- 2.95924e-39 + -6.63424e-39 = -3.675e-39
	(b"10000000010111010011111111010010", b"00000000000000000000000000000000"),
	(b"10000000011100010011010101001110", b"10000000110011100111010100100000"), -- -8.5636e-39 + -1.03965e-38 = -1.89601e-38
	(b"10000000011111100011101001101000", b"00000000000000000000000000000000"),
	(b"00000000001100110000001010101010", b"10000000010010110011011110111110"), -- -1.15922e-38 + 4.68457e-39 = -6.90766e-39
	(b"00000000010010111111110101001111", b"00000000000000000000000000000000"),
	(b"10000000010000000001011011101111", b"00000000000010111110011001100000"), -- 6.97853e-39 + -5.8857e-39 = 1.09283e-39
	(b"00000000010011010100101100110000", b"00000000000000000000000000000000"),
	(b"10000000000101000011001000111001", b"00000000001110010001100011110111"), -- 7.09831e-39 + -1.85473e-39 = 5.24358e-39
	(b"00000000010001100010000110001110", b"00000000000000000000000000000000"),
	(b"10000000000111011000100000101000", b"00000000001010001001100101100110"), -- 6.44052e-39 + -2.71207e-39 = 3.72845e-39
	(b"00000000000100001111000100001000", b"00000000000000000000000000000000"),
	(b"10000000000010011111000001011010", b"00000000000001110000000010101110"), -- 1.55583e-39 + -9.12741e-40 = 6.43092e-40
	(b"00000000010101010011010010100100", b"00000000000000000000000000000000"),
	(b"10000000000010101111111101100011", b"00000000010010100011010101000001"), -- 7.8249e-39 + -1.00997e-39 = 6.81493e-39
	(b"10000000010110100011110111100110", b"00000000000000000000000000000000"),
	(b"10000000001011011011001001000101", b"10000000100001111111000000101011"), -- -8.2874e-39 + -4.19655e-39 = -1.24839e-38
	(b"00000000010100001001111011111101", b"00000000000000000000000000000000"),
	(b"10000000011011001111110111001000", b"10000000000111000101111011001011"), -- 7.40387e-39 + -1.00093e-38 = -2.6054e-39
	(b"10000000011101101110000000011001", b"00000000000000000000000000000000"),
	(b"00000000010010011001100000100110", b"10000000001011010100011111110011"), -- -1.0917e-38 + 6.75857e-39 = -4.15841e-39
	(b"00000000000010011001010101101101", b"00000000000000000000000000000000"),
	(b"10000000001010010011101000010100", b"10000000000111111010010010100111"), -- 8.80123e-40 + -3.78609e-39 = -2.90597e-39
	(b"10000000011110101111111010001111", b"00000000000000000000000000000000"),
	(b"10000000001011101111001000010100", b"10000000101010011111000010100011"), -- -1.12952e-38 + -4.31127e-39 = -1.56065e-38
	(b"00000000010110100001010010100001", b"00000000000000000000000000000000"),
	(b"10000000000110001000000101100001", b"00000000010000011001001101000000"), -- 8.27259e-39 + -2.25046e-39 = 6.02213e-39
	(b"10000000000111101111000101011100", b"00000000000000000000000000000000"),
	(b"00000000011001010100111000100101", b"00000000010001100101110011001001"), -- -2.84165e-39 + 9.30342e-39 = 6.46177e-39
	(b"00000000001111101101101011110111", b"00000000000000000000000000000000"),
	(b"10000000011001100011011000001101", b"10000000001001110101101100010110"), -- 5.77235e-39 + -9.38661e-39 = -3.61426e-39
	(b"00000000010000001101000101000111", b"00000000000000000000000000000000"),
	(b"10000000000111001100100010001100", b"00000000001001000000100010111011"), -- 5.95255e-39 + -2.64334e-39 = 3.30921e-39
	(b"10000000001100100111010001000110", b"00000000000000000000000000000000"),
	(b"10000000001011011001110010001001", b"10000000011000000001000011001111"), -- -4.63349e-39 + -4.18875e-39 = -8.82224e-39
	(b"10000000000010111001010000111000", b"00000000000000000000000000000000"),
	(b"10000000001110001011101011010100", b"10000000010001000100111100001100"), -- -1.06336e-39 + -5.20981e-39 = -6.27317e-39
	(b"10000000011110111010001001100000", b"00000000000000000000000000000000"),
	(b"10000000011111110101001011010001", b"10000000111110101111010100110001"), -- -1.1354e-38 + -1.16928e-38 = -2.30468e-38
	(b"00000000011101010010010100000101", b"00000000000000000000000000000000"),
	(b"10000000000011000110001111101110", b"00000000011010001100000100010111"), -- 1.0758e-38 + -1.13787e-39 = 9.62016e-39
	(b"10000000001100111011111101000000", b"00000000000000000000000000000000"),
	(b"10000000001100010101101011000101", b"10000000011001010001101000000101"), -- -4.75222e-39 + -4.5325e-39 = -9.28472e-39
	(b"10000000000011110101100111000100", b"00000000000000000000000000000000"),
	(b"00000000010111110111110111101010", b"00000000010100000010010000100110"), -- -1.40973e-39 + 8.76954e-39 = 7.35981e-39
	(b"00000000000000110101001000000000", b"00000000000000000000000000000000"),
	(b"10000000000101000101000111101101", b"10000000000100001111111111101101"), -- 3.04923e-40 + -1.8661e-39 = -1.56118e-39
	(b"10000000011101001101011001110011", b"00000000000000000000000000000000"),
	(b"10000000011101110000000001000100", b"10000000111010111101011010110111"), -- -1.07298e-38 + -1.09285e-38 = -2.16584e-38
	(b"10000000011010001110110110111101", b"00000000000000000000000000000000"),
	(b"00000000010100011010000011101010", b"10000000000101110100110011010011"), -- -9.63618e-39 + 7.4964e-39 = -2.13978e-39
	(b"10000000000000001110000010100101", b"00000000000000000000000000000000"),
	(b"10000000000110111001100110010000", b"10000000000111000111101000110101"), -- -8.05873e-41 + -2.53465e-39 = -2.61523e-39
	(b"10000000010110101000100010101110", b"00000000000000000000000000000000"),
	(b"10000000000111011011100111110100", b"10000000011110000100001010100010"), -- -8.31423e-39 + -2.72994e-39 = -1.10442e-38
	(b"10000000010110010001000011110111", b"00000000000000000000000000000000"),
	(b"00000000010111111101001110101001", b"00000000000001101100001010110010"), -- -8.17944e-39 + 8.8003e-39 = 6.20856e-40
	(b"00000000011110000110100101001111", b"00000000000000000000000000000000"),
	(b"10000000001011010101100001001011", b"00000000010010110001000100000100"), -- 1.1058e-38 + -4.16427e-39 = 6.89377e-39
	(b"10000000001001001101100010100111", b"00000000000000000000000000000000"),
	(b"10000000010010011100110010010001", b"10000000011011101010010100111000"), -- -3.3838e-39 + -6.77738e-39 = -1.01612e-38
	(b"10000000010000011100111111001000", b"00000000000000000000000000000000"),
	(b"10000000010111001000100110100011", b"10000000100111100101100101101011"), -- -6.04385e-39 + -8.49824e-39 = -1.45421e-38
	(b"10000000011000101011110111001011", b"00000000000000000000000000000000"),
	(b"10000000000111010000110100100111", b"10000000011111111100101011110010"), -- -9.06796e-39 + -2.66795e-39 = -1.17359e-38
	(b"00000000011110101001001110111110", b"00000000000000000000000000000000"),
	(b"10000000010101001111010110100101", b"00000000001001011001111000011001"), -- 1.12569e-38 + -7.8023e-39 = 3.45463e-39
	(b"00000000010001011000011001111111", b"00000000000000000000000000000000"),
	(b"10000000010010011111110000010100", b"10000000000001000111010110010101"), -- 6.3849e-39 + -6.79442e-39 = -4.09522e-40
	(b"00000000000010111001001101001100", b"00000000000000000000000000000000"),
	(b"10000000000110101010101001011111", b"10000000000011110001011100010011"), -- 1.06303e-39 + -2.44884e-39 = -1.38581e-39
	(b"10000000001000111111100111110001", b"00000000000000000000000000000000"),
	(b"10000000000001011000101101100111", b"10000000001010011000010101011000"), -- -3.3039e-39 + -5.09186e-40 = -3.81309e-39
	(b"00000000001111110101111010110111", b"00000000000000000000000000000000"),
	(b"10000000000001110011101100010010", b"00000000001110000010001110100101"), -- 5.81961e-39 + -6.64039e-40 = 5.15557e-39
	(b"00000000000001110101100101010110", b"00000000000000000000000000000000"),
	(b"10000000000111010000001111000110", b"10000000000101011010101001110000"), -- 6.74896e-40 + -2.66458e-39 = -1.98969e-39
	(b"10000000010011101010011111001101", b"00000000000000000000000000000000"),
	(b"00000000001011011011000100000010", b"10000000001000001111011011001011"), -- -7.22336e-39 + 4.1961e-39 = -3.02727e-39
	(b"10000000010001010101100000110111", b"00000000000000000000000000000000"),
	(b"00000000001110011000100101000111", b"10000000000010111100111011110000"), -- -6.36829e-39 + 5.28387e-39 = -1.08443e-39
	(b"00000000001110001110000110101101", b"00000000000000000000000000000000"),
	(b"10000000001100010010010110001110", b"00000000000001111011110000011111"), -- 5.22375e-39 + -4.51341e-39 = 7.10334e-40
	(b"10000000011111110110110100010001", b"00000000000000000000000000000000"),
	(b"10000000010101011100111000111001", b"10000000110101010011101101001010"), -- -1.17022e-38 + -7.88e-39 = -1.95822e-38
	(b"00000000001000100000101100101010", b"00000000000000000000000000000000"),
	(b"00000000000011100010001100110010", b"00000000001100000010111001011100"), -- 3.12641e-39 + 1.29832e-39 = 4.42473e-39
	(b"00000000000001011110000110011010", b"00000000000000000000000000000000"),
	(b"00000000001111011001111010101011", b"00000000010000111000000001000101"), -- 5.40108e-40 + 5.65888e-39 = 6.19899e-39
	(b"10000000011010000100001111001110", b"00000000000000000000000000000000"),
	(b"10000000010001110000001101100000", b"10000000101011110100011100101110"), -- -9.57522e-39 + -6.52153e-39 = -1.60967e-38
	(b"00000000000010110010001100111001", b"00000000000000000000000000000000"),
	(b"10000000001000001000111101100101", b"10000000000101010110110000101100"), -- 1.02283e-39 + -2.99018e-39 = -1.96735e-39
	(b"00000000011100101111101110001100", b"00000000000000000000000000000000"),
	(b"10000000010110110111011111000001", b"00000000000101111000001111001011"), -- 1.05595e-38 + -8.39999e-39 = 2.15949e-39
	(b"10000000010111100010000101001111", b"00000000000000000000000000000000"),
	(b"00000000011011111110111101010100", b"00000000000100011100111000000101"), -- -8.64449e-39 + 1.02796e-38 = 1.63511e-39
	(b"00000000000011010010001111010001", b"00000000000000000000000000000000"),
	(b"10000000010101001010000100101101", b"10000000010001110111110101011100"), -- 1.20671e-39 + -7.772e-39 = -6.56529e-39
	(b"10000000010000010100110000111011", b"00000000000000000000000000000000"),
	(b"10000000010010100000001011000010", b"10000000100010110100111011111101"), -- -5.99665e-39 + -6.79682e-39 = -1.27935e-38
	(b"10000000000010010110001000100010", b"00000000000000000000000000000000"),
	(b"10000000000100111000100010100001", b"10000000000111001110101011000011"), -- -8.61723e-40 + -1.79389e-39 = -2.65561e-39
	(b"10000000010101000101100001000100", b"00000000000000000000000000000000"),
	(b"00000000000100011001101100011011", b"10000000010000101011110100101001"), -- -7.74585e-39 + 1.61684e-39 = -6.129e-39
	(b"10000000011010011001001010000011", b"00000000000000000000000000000000"),
	(b"00000000011000101001101011110010", b"10000000000001101111011110010001"), -- -9.69529e-39 + 9.05546e-39 = -6.39823e-40
	(b"10000000011011110111101001000010", b"00000000000000000000000000000000"),
	(b"00000000010001010010010001110001", b"10000000001010100101010111010001"), -- -1.02376e-38 + 6.34972e-39 = -3.88788e-39
	(b"00000000010000111101001111011011", b"00000000000000000000000000000000"),
	(b"10000000001001001111101001001100", b"00000000000111101101100110001111"), -- 6.22898e-39 + -3.39587e-39 = 2.83311e-39
	(b"10000000001111101110010011001101", b"00000000000000000000000000000000"),
	(b"10000000011100000100000000111110", b"10000000101011110010010100001011"), -- -5.77588e-39 + -1.03086e-38 = -1.60845e-38
	(b"00000000000101101111111111001011", b"00000000000000000000000000000000"),
	(b"00000000001111001000111111110100", b"00000000010100111000111110111111"), -- 2.11214e-39 + 5.56177e-39 = 7.67391e-39
	(b"10000000011111101111000001100111", b"00000000000000000000000000000000"),
	(b"00000000000000010001110001010111", b"10000000011111011101010000010000"), -- -1.16575e-38 + 1.02002e-40 = -1.15555e-38
	(b"10000000011000000000110101100100", b"00000000000000000000000000000000"),
	(b"00000000000010001111111000100010", b"10000000010101110000111101000010"), -- -8.82101e-39 + 8.2585e-40 = -7.99516e-39
	(b"00000000000000001000111101010010", b"00000000000000000000000000000000"),
	(b"10000000010001101101010000111101", b"10000000010001100100010011101011"), -- 5.14136e-41 + -6.50462e-39 = -6.45321e-39
	(b"10000000001000111001100111000010", b"00000000000000000000000000000000"),
	(b"10000000011111100010101111011011", b"10000000101000011100010110011101"), -- -3.2694e-39 + -1.1587e-38 = -1.48564e-38
	(b"10000000001101110101100111111000", b"00000000000000000000000000000000"),
	(b"10000000011010111110111110010011", b"10000000101000110100100110001011"), -- -5.08323e-39 + -9.91234e-39 = -1.49956e-38
	(b"10000000011101111011111001111100", b"00000000000000000000000000000000"),
	(b"00000000010000010001111100000010", b"10000000001101101001111101111010"), -- -1.09968e-38 + 5.98043e-39 = -5.01633e-39
	(b"10000000010111000111010011001101", b"00000000000000000000000000000000"),
	(b"10000000010100010101110100100000", b"10000000101011011101000111101101"), -- -8.49077e-39 + -7.47208e-39 = -1.59628e-38
	(b"10000000000101110011100110000011", b"00000000000000000000000000000000"),
	(b"00000000010111000011001010010110", b"00000000010001001111100100010011"), -- -2.13285e-39 + 8.46701e-39 = 6.33416e-39
	(b"00000000011010011100101111011011", b"00000000000000000000000000000000"),
	(b"10000000011100110010010101101011", b"10000000000010010101100110010000"), -- 9.71586e-39 + -1.05745e-38 = -8.58648e-40
	(b"10000000010101000011110100110010", b"00000000000000000000000000000000"),
	(b"10000000001011010101000011000101", b"10000000100000011000110111110111"), -- -7.73613e-39 + -4.16157e-39 = -1.18977e-38
	(b"00000000000000010000110100101100", b"00000000000000000000000000000000"),
	(b"10000000001011010011011001001011", b"10000000001011000010100100011111"), -- 9.65607e-41 + -4.15207e-39 = -4.05551e-39
	(b"00000000010110011001110110000010", b"00000000000000000000000000000000"),
	(b"10000000001001101010110010110010", b"00000000001100101111000011010000"), -- 8.22986e-39 + -3.5517e-39 = 4.67816e-39
	(b"10000000011001101100110001011110", b"00000000000000000000000000000000"),
	(b"00000000000111000011011100001010", b"10000000010010101001010101010100"), -- -9.44053e-39 + 2.59114e-39 = -6.8494e-39
	(b"10000000000001011100010001101011", b"00000000000000000000000000000000"),
	(b"00000000010010100001111100001011", b"00000000010001000101101010100000"), -- -5.29639e-40 + 6.80696e-39 = 6.27732e-39
	(b"10000000010110101010010010010010", b"00000000000000000000000000000000"),
	(b"00000000010000000000010010100011", b"10000000000110101001111111101111"), -- -8.32423e-39 + 5.87914e-39 = -2.4451e-39
	(b"00000000011101111011101001001011", b"00000000000000000000000000000000"),
	(b"00000000000101010001011111110001", b"00000000100011001101001000111100"), -- 1.09953e-38 + 1.93713e-39 = 1.29324e-38
	(b"10000000010011101100011111001101", b"00000000000000000000000000000000"),
	(b"00000000010101010011101101010011", b"00000000000001100111001110000110"), -- -7.23484e-39 + 7.8273e-39 = 5.92455e-40
	(b"10000000010111101011101110100100", b"00000000000000000000000000000000"),
	(b"10000000000110010110000010011001", b"10000000011110000001110000111101"), -- -8.69985e-39 + -2.33054e-39 = -1.10304e-38
	(b"10000000001011100110000111100101", b"00000000000000000000000000000000"),
	(b"10000000011111010000001001011001", b"10000000101010110110010000111110"), -- -4.25955e-39 + -1.14803e-38 = -1.57398e-38
	(b"00000000010101001111010010001000", b"00000000000000000000000000000000"),
	(b"00000000001110011000000011001001", b"00000000100011100111010101010001"), -- 7.8019e-39 + 5.28082e-39 = 1.30827e-38
	(b"00000000011001010010001110010110", b"00000000000000000000000000000000"),
	(b"10000000011010011001100000011101", b"10000000000001000111010010000111"), -- 9.28815e-39 + -9.6973e-39 = -4.09144e-40
	(b"00000000010100111001110011000010", b"00000000000000000000000000000000"),
	(b"10000000001100001011011000101011", b"00000000001000101110011010010111"), -- 7.67858e-39 + -4.47345e-39 = 3.20513e-39
	(b"10000000011001001101011111111100", b"00000000000000000000000000000000"),
	(b"10000000000100000111111110100011", b"10000000011101010101011110011111"), -- -9.26103e-39 + -1.51516e-39 = -1.07762e-38
	(b"10000000001100100110000011010110", b"00000000000000000000000000000000"),
	(b"00000000001100000001011010100011", b"10000000000000100100101000110011"), -- -4.62651e-39 + 4.41622e-39 = -2.10289e-40
	(b"00000000000011101010100011001111", b"00000000000000000000000000000000"),
	(b"00000000001010101001111000101011", b"00000000001110010100011011111010"), -- 1.34625e-39 + 3.91383e-39 = 5.26008e-39
	(b"10000000010100011111111010000010", b"00000000000000000000000000000000"),
	(b"10000000011010110111100110101001", b"10000000101111010111100000101011"), -- -7.52998e-39 + -9.87004e-39 = -1.74e-38
	(b"00000000011111000101000010111001", b"00000000000000000000000000000000"),
	(b"00000000011011010111000011001111", b"00000000111010011100000110001000"), -- 1.14166e-38 + 1.00505e-38 = 2.14671e-38
	(b"00000000010000110110110111100101", b"00000000000000000000000000000000"),
	(b"10000000010000110001001101000101", b"00000000000000000101101010100000"), -- 6.1924e-39 + -6.15989e-39 = 3.25101e-41
	(b"00000000011111111010110000001001", b"00000000000000000000000000000000"),
	(b"00000000010011111110001100100111", b"00000000110011111000111100110000"), -- 1.17248e-38 + 7.33649e-39 = 1.90613e-38
	(b"10000000010000000110100000110101", b"00000000000000000000000000000000"),
	(b"10000000011110011110001001001101", b"10000000101110100100101010000010"), -- -5.91485e-39 + -1.11933e-38 = -1.71081e-38
	(b"10000000000001111011101101001111", b"00000000000000000000000000000000"),
	(b"10000000001110011000000110001101", b"10000000010000010011110011011100"), -- -7.10042e-40 + -5.2811e-39 = -5.99114e-39
	(b"00000000011110110100000101110011", b"00000000000000000000000000000000"),
	(b"00000000010010011101001001001100", b"00000000110001010001001110111111"), -- 1.13192e-38 + 6.77943e-39 = 1.80987e-38
	(b"10000000001001011000110110000001", b"00000000000000000000000000000000"),
	(b"10000000001010000011111000101101", b"10000000010011011100101110101110"), -- -3.44868e-39 + -3.69572e-39 = -7.1444e-39
	(b"10000000001111011000110100011111", b"00000000000000000000000000000000"),
	(b"00000000001111101111101110000011", b"00000000000000010110111001100100"), -- -5.65259e-39 + 5.78403e-39 = 1.31436e-40
	(b"00000000001110100111101101110000", b"00000000000000000000000000000000"),
	(b"00000000011011101110110000000100", b"00000000101010010110011101110100"), -- 5.37074e-39 + 1.01866e-38 = 1.55573e-38
	(b"00000000011011100001011110101001", b"00000000000000000000000000000000"),
	(b"00000000001011001001100011101011", b"00000000100110101011000010010100"), -- 1.01104e-38 + 4.09562e-39 = 1.4206e-38
	(b"10000000001110000111000001111111", b"00000000000000000000000000000000"),
	(b"10000000001011001001100110111010", b"10000000011001010000101000111001"), -- -5.18314e-39 + -4.09591e-39 = -9.27905e-39
	(b"10000000001100010100000000100101", b"00000000000000000000000000000000"),
	(b"00000000001010000100100110001001", b"10000000000010001111011010011100"), -- -4.52295e-39 + 3.6998e-39 = -8.23151e-40
	(b"10000000010111011001010001101011", b"00000000000000000000000000000000"),
	(b"00000000010110000110011000111010", b"10000000000001010010111000110001"), -- -8.59394e-39 + 8.1182e-39 = -4.75748e-40
	(b"10000000000101000110111101100111", b"00000000000000000000000000000000"),
	(b"00000000001010111011010000000010", b"00000000000101110100010010011011"), -- -1.87667e-39 + 4.0135e-39 = 2.13683e-39
	(b"10000000001110000000110010000100", b"00000000000000000000000000000000"),
	(b"10000000011111111100001011110001", b"10000000101101111100111101110101"), -- -5.14728e-39 + -1.1733e-38 = -1.68803e-38
	(b"00000000010110101111011101111000", b"00000000000000000000000000000000"),
	(b"10000000010101111101010110111001", b"00000000000000110010000110111111"), -- 8.35397e-39 + -8.06636e-39 = 2.87612e-40
	(b"10000000010101111010111001000010", b"00000000000000000000000000000000"),
	(b"00000000001010000000101001010100", b"10000000001011111010001111101110"), -- -8.0522e-39 + 3.67712e-39 = -4.37508e-39
	(b"10000000000111110011101111111010", b"00000000000000000000000000000000"),
	(b"10000000011010010101101000010000", b"10000000100010001001011000001010"), -- -2.86842e-39 + -9.67504e-39 = -1.25435e-38
	(b"00000000001101010110101010111110", b"00000000000000000000000000000000"),
	(b"00000000001111100100110001101010", b"00000000011100111011011100101000"), -- 4.90557e-39 + 5.72121e-39 = 1.06268e-38
	(b"00000000011111101010001011111000", b"00000000000000000000000000000000"),
	(b"10000000011011111111000111000100", b"00000000000011101011000100110100"), -- 1.16297e-38 + -1.02805e-38 = 1.34927e-39
	(b"10000000010010001000111010010110", b"00000000000000000000000000000000"),
	(b"00000000011111011001100011010101", b"00000000001101010000101000111111"), -- -6.66331e-39 + 1.15343e-38 = 4.87096e-39
	(b"00000000011011011101100111101011", b"00000000000000000000000000000000"),
	(b"00000000011001010100010110110001", b"00000000110100110001111110011100"), -- 1.00882e-38 + 9.30039e-39 = 1.93886e-38
	(b"10000000000011111111101011001100", b"00000000000000000000000000000000"),
	(b"00000000001101111011001111010110", b"00000000001001111011100100001010"), -- -1.4675e-39 + 5.11547e-39 = 3.64796e-39
	(b"00000000000100001101001001000101", b"00000000000000000000000000000000"),
	(b"00000000001111000100110001101000", b"00000000010011010001111010101101"), -- 1.5448e-39 + 5.53754e-39 = 7.08234e-39
	(b"00000000001100110110100000011111", b"00000000000000000000000000000000"),
	(b"00000000001011000111010101010000", b"00000000010111111101110101101111"), -- 4.72096e-39 + 4.08285e-39 = 8.80381e-39
	(b"10000000001111111000111000100011", b"00000000000000000000000000000000"),
	(b"00000000010001000100111010101111", b"00000000000001001100000010001100"), -- -5.83663e-39 + 6.27304e-39 = 4.36415e-40
	(b"00000000000001111111011011000111", b"00000000000000000000000000000000"),
	(b"10000000000101000001001101011010", b"10000000000011000001110010010011"), -- 7.31376e-40 + -1.84365e-39 = -1.11228e-39
	(b"10000000010010001010111101010000", b"00000000000000000000000000000000"),
	(b"00000000001111100110100101011000", b"10000000000010100100010111111000"), -- -6.67505e-39 + 5.73159e-39 = -9.43455e-40
	(b"00000000000111110000100100000011", b"00000000000000000000000000000000"),
	(b"00000000001010010110101100101001", b"00000000010010000111010000101100"), -- 2.85013e-39 + 3.8037e-39 = 6.65383e-39
	(b"10000000010110011000011011101101", b"00000000000000000000000000000000"),
	(b"10000000001001010100001111011011", b"10000000011111101100101011001000"), -- -8.22176e-39 + -3.42226e-39 = -1.1644e-38
	(b"10000000011011001011011101101010", b"00000000000000000000000000000000"),
	(b"10000000000010010101110001101011", b"10000000011101100001001111010101"), -- -9.98403e-39 + -8.59673e-40 = -1.08437e-38
	(b"00000000011011100011000011010010", b"00000000000000000000000000000000"),
	(b"10000000011001111111111101001000", b"00000000000001100011000110001010"), -- 1.01194e-38 + -9.55063e-39 = 5.68784e-40
	(b"10000000010111101110001100111110", b"00000000000000000000000000000000"),
	(b"00000000001011000000100000111110", b"10000000001100101101101100000000"), -- -8.71406e-39 + 4.04372e-39 = -4.67034e-39
	(b"10000000010011001101111001000010", b"00000000000000000000000000000000"),
	(b"00000000000000110111000110101100", b"10000000010010010110110010010110"), -- -7.05923e-39 + 3.16284e-40 = -6.74294e-39
	(b"10000000001100101000101011001111", b"00000000000000000000000000000000"),
	(b"00000000011110010001101101110111", b"00000000010001101001000010101000"), -- -4.64157e-39 + 1.11219e-38 = 6.48038e-39
	(b"00000000010010000110011100111000", b"00000000000000000000000000000000"),
	(b"10000000001000100100111111000000", b"00000000001001100001011101111000"), -- 6.64918e-39 + -3.15102e-39 = 3.49817e-39
	(b"00000000000001101101110101111011", b"00000000000000000000000000000000"),
	(b"00000000010100011110101010101001", b"00000000010110001100100000100100"), -- 6.30465e-40 + 7.52286e-39 = 8.15332e-39
	(b"00000000001101011000010000001011", b"00000000000000000000000000000000"),
	(b"10000000011101111101011101011111", b"10000000010000100101001101010100"), -- 4.91465e-39 + -1.10057e-38 = -6.09104e-39
	(b"10000000001101100100111000101110", b"00000000000000000000000000000000"),
	(b"10000000010100111011011111001001", b"10000000100010100000010111110111"), -- -4.98716e-39 + -7.68828e-39 = -1.26754e-38
	(b"00000000000000111010101001001001", b"00000000000000000000000000000000"),
	(b"10000000010001100011010010000010", b"10000000010000101000101000111001"), -- 3.36593e-40 + -6.44732e-39 = -6.11073e-39
	(b"10000000001101011001110001000000", b"00000000000000000000000000000000"),
	(b"10000000010100111101101111010000", b"10000000100010010111100000010000"), -- -4.92333e-39 + -7.7012e-39 = -1.26245e-38
	(b"00000000011110111111110000011111", b"00000000000000000000000000000000"),
	(b"10000000010000100101110111000000", b"00000000001110011001111001011111"), -- 1.13862e-38 + -6.09477e-39 = 5.29144e-39
	(b"10000000011000100101010100110111", b"00000000000000000000000000000000"),
	(b"10000000011011110111111010010000", b"10000000110100011101001111000111"), -- -9.03045e-39 + -1.02391e-38 = -1.92696e-38
	(b"00000000011000010110111111100010", b"00000000000000000000000000000000"),
	(b"10000000010110111100101110000100", b"00000000000001011010010001011110"), -- 8.94818e-39 + -8.43004e-39 = 5.18141e-40
	(b"00000000011011000011110000001110", b"00000000000000000000000000000000"),
	(b"00000000011011011110010000111101", b"00000000110110100010000001001011"), -- 9.93978e-39 + 1.00919e-38 = 2.00317e-38
	(b"10000000011001010001010000011011", b"00000000000000000000000000000000"),
	(b"00000000010001110101001000011111", b"10000000000111011100000111111100"), -- -9.2826e-39 + 6.54978e-39 = -2.73282e-39
	(b"10000000000110010011011110100000", b"00000000000000000000000000000000"),
	(b"10000000001001001000110000001101", b"10000000001111011100001110101101"), -- -2.31584e-39 + -3.35632e-39 = -5.67216e-39
	(b"00000000010011000101010000100101", b"00000000000000000000000000000000"),
	(b"00000000001011100101101000101000", b"00000000011110101010111001001101"), -- 7.00968e-39 + 4.25677e-39 = 1.12665e-38
	(b"00000000000110010111011111111101", b"00000000000000000000000000000000"),
	(b"10000000000010100001101011010111", b"00000000000011110101110100100110"), -- 2.33893e-39 + -9.27983e-40 = 1.41095e-39
	(b"10000000001001011001000100101101", b"00000000000000000000000000000000"),
	(b"00000000010100110010001110110100", b"00000000001011011001001010000111"), -- -3.44999e-39 + 7.63515e-39 = 4.18516e-39
	(b"00000000010101001010101001101000", b"00000000000000000000000000000000"),
	(b"00000000001000000111111111100111", b"00000000011101010010101001001111"), -- 7.77531e-39 + 2.98462e-39 = 1.07599e-38
	(b"00000000010100011001001010100010", b"00000000000000000000000000000000"),
	(b"10000000011001110101101001101011", b"10000000000101011100011111001001"), -- 7.49128e-39 + -9.49149e-39 = -2.00021e-39
	(b"10000000010000100110101010000100", b"00000000000000000000000000000000"),
	(b"00000000001011111101011110010011", b"10000000000100101001001011110001"), -- -6.09935e-39 + 4.3936e-39 = -1.70575e-39
	(b"00000000010101001111000111010100", b"00000000000000000000000000000000"),
	(b"10000000001100100010100101111000", b"00000000001000101100100001011100"), -- 7.80093e-39 + -4.60665e-39 = 3.19428e-39
	(b"00000000001110011101111010010001", b"00000000000000000000000000000000"),
	(b"10000000011111001011001001111110", b"10000000010000101101001111101101"), -- 5.31447e-39 + -1.14516e-38 = -6.13717e-39
	(b"00000000011000100010000001010011", b"00000000000000000000000000000000"),
	(b"10000000010100111101000110100101", b"00000000000011100100111010101110"), -- 9.01147e-39 + -7.69755e-39 = 1.31392e-39
	(b"00000000001001000100101111111011", b"00000000000000000000000000000000"),
	(b"00000000010100001011011100000001", b"00000000011101010000001011111100"), -- 3.33333e-39 + 7.41249e-39 = 1.07458e-38
	(b"00000000001101010010011110011100", b"00000000000000000000000000000000"),
	(b"10000000010110011010110000101000", b"10000000001001001000010010001100"), -- 4.88149e-39 + -8.23512e-39 = -3.35363e-39
	(b"00000000001101010101011010111101", b"00000000000000000000000000000000"),
	(b"10000000000110111010111010001011", b"00000000000110011010100000110010"), -- 4.8984e-39 + -2.54217e-39 = 2.35622e-39
	(b"00000000000110111001100100011011", b"00000000000000000000000000000000"),
	(b"10000000011110100101110100001100", b"10000000010111101100001111110001"), -- 2.53448e-39 + -1.12373e-38 = -8.70283e-39
	(b"10000000011100001000001111001101", b"00000000000000000000000000000000"),
	(b"00000000011010000111111011111101", b"10000000000010000000010011010000"), -- -1.03329e-38 + 9.59645e-39 = -7.3641e-40
	(b"00000000001010010100101010100011", b"00000000000000000000000000000000"),
	(b"10000000010110111110100101001110", b"10000000001100101001111010101011"), -- 3.79203e-39 + -8.44072e-39 = -4.64869e-39
	(b"00000000011101000110010100011000", b"00000000000000000000000000000000"),
	(b"10000000011110100000110110010010", b"10000000000001011010100001111010"), -- 1.06892e-38 + -1.12088e-38 = -5.19615e-40
	(b"10000000011100001001011011101111", b"00000000000000000000000000000000"),
	(b"10000000010111010101100110000111", b"10000000110011011111000001110110"), -- -1.03397e-38 + -8.57282e-39 = -1.89125e-38
	(b"10000000011000010000001110110001", b"00000000000000000000000000000000"),
	(b"10000000001000010110000100110011", b"10000000100000100110010011100100"), -- -8.90937e-39 + -3.06544e-39 = -1.19748e-38
	(b"00000000001010000001010011101001", b"00000000000000000000000000000000"),
	(b"10000000001110001101100010001110", b"10000000000100001100001110100101"), -- 3.68092e-39 + -5.22047e-39 = -1.53955e-39
	(b"00000000011001011111011001101011", b"00000000000000000000000000000000"),
	(b"10000000011011001010000011100001", b"10000000000001101010101001110110"), -- 9.36378e-39 + -9.97595e-39 = -6.12163e-40
	(b"00000000011101001110010101011001", b"00000000000000000000000000000000"),
	(b"10000000001111100010111011000010", b"00000000001101101011011010010111"), -- 1.07352e-38 + -5.71057e-39 = 5.02462e-39
	(b"10000000011110001011011010011001", b"00000000000000000000000000000000"),
	(b"10000000011101101011101000100101", b"10000000111011110111000010111110"), -- -1.10858e-38 + -1.09034e-38 = -2.19891e-38
	(b"10000000010111111101101110111111", b"00000000000000000000000000000000"),
	(b"00000000010011110111001010100111", b"10000000000100000110100100011000"), -- -8.8032e-39 + 7.29613e-39 = -1.50707e-39
	(b"10000000001110011010001000111010", b"00000000000000000000000000000000"),
	(b"10000000000101111001000111001110", b"10000000010100010011010000001000"), -- -5.29282e-39 + -2.16452e-39 = -7.45734e-39
	(b"00000000010111100010001000111000", b"00000000000000000000000000000000"),
	(b"10000000011110001111011011101101", b"10000000000110101101010010110101"), -- 8.64481e-39 + -1.11088e-38 = -2.46403e-39
	(b"10000000011111000111011001010000", b"00000000000000000000000000000000"),
	(b"00000000010011011111110111111010", b"10000000001011100111100001010110"), -- -1.143e-38 + 7.16244e-39 = -4.2676e-39
	(b"10000000011000001000001100001101", b"00000000000000000000000000000000"),
	(b"00000000010100010111011101110100", b"10000000000011110000101110011001"), -- -8.86322e-39 + 7.48153e-39 = -1.38169e-39
	(b"00000000000100111010001100111000", b"00000000000000000000000000000000"),
	(b"10000000001010110101100011011101", b"10000000000101111011010110100101"), -- 1.80343e-39 + -3.9808e-39 = -2.17738e-39
	(b"00000000010011010000001110010101", b"00000000000000000000000000000000"),
	(b"00000000010101111010000111010010", b"00000000101001001010010101100111"), -- 7.07262e-39 + 8.04774e-39 = 1.51204e-38
	(b"00000000001010001110011111010100", b"00000000000000000000000000000000"),
	(b"10000000010111001101110100011111", b"10000000001100111111010101001011"), -- 3.75658e-39 + -8.52819e-39 = -4.7716e-39
	(b"10000000000110110101101100110001", b"00000000000000000000000000000000"),
	(b"00000000010001000111111010101101", b"00000000001010010010001101111100"), -- -2.51227e-39 + 6.29026e-39 = 3.77798e-39
	(b"00000000001011110011110100001011", b"00000000000000000000000000000000"),
	(b"10000000011011111101111110111110", b"10000000010000001010001010110011"), -- 4.33817e-39 + -1.0274e-38 = -5.93584e-39
	(b"00000000011110001001111011000011", b"00000000000000000000000000000000"),
	(b"00000000000000010011000011110111", b"00000000011110011100111110111010"), -- 1.10772e-38 + 1.09401e-40 = 1.11866e-38
	(b"10000000000010100111000010000111", b"00000000000000000000000000000000"),
	(b"10000000011110100100001111110111", b"10000000100001001011010001111110"), -- -9.58722e-40 + -1.12283e-38 = -1.2187e-38
	(b"00000000011011001110011011011011", b"00000000000000000000000000000000"),
	(b"00000000000111110010110110101100", b"00000000100011000001010010000111"), -- 1.0001e-38 + 2.86328e-39 = 1.28643e-38
	(b"10000000010000011000000001001100", b"00000000000000000000000000000000"),
	(b"10000000010110100101100100001001", b"10000000100110111101100101010101"), -- -6.01533e-39 + -8.29713e-39 = -1.43125e-38
	(b"00000000010010101000001111100010", b"00000000000000000000000000000000"),
	(b"10000000011111110111101011111110", b"10000000001101001111011100011100"), -- 6.84314e-39 + -1.17072e-38 = -4.86409e-39
	(b"00000000000010000110000010000101", b"00000000000000000000000000000000"),
	(b"00000000001101100101011101101111", b"00000000001111101011011111110100"), -- 7.69309e-40 + 4.99048e-39 = 5.75979e-39
	(b"10000000001110000100010100001110", b"00000000000000000000000000000000"),
	(b"00000000000011100001100011000110", b"10000000001010100010110001001000"), -- -5.16756e-39 + 1.29458e-39 = -3.87298e-39
	(b"10000000010110010111110101001111", b"00000000000000000000000000000000"),
	(b"00000000000000101001101101000100", b"10000000010101101110001000001011"), -- -8.21831e-39 + 2.3937e-40 = -7.97894e-39
	(b"00000000001111000110111101100100", b"00000000000000000000000000000000"),
	(b"00000000011010011001001101111101", b"00000000101001100000001011100001"), -- 5.55009e-39 + 9.69564e-39 = 1.52457e-38
	(b"10000000000110010010011011000010", b"00000000000000000000000000000000"),
	(b"10000000001001110000110111001011", b"10000000010000000011010010001101"), -- -2.30979e-39 + -3.58653e-39 = -5.89632e-39
	(b"00000000001111010000000011010111", b"00000000000000000000000000000000"),
	(b"10000000010001010110001010001100", b"10000000000010000110000110110101"), -- 5.60227e-39 + -6.372e-39 = -7.69735e-40
	(b"10000000011101001001011010010100", b"00000000000000000000000000000000"),
	(b"10000000001011110101010111001000", b"10000000101000111110110001011100"), -- -1.07069e-38 + -4.34704e-39 = -1.5054e-38
	(b"10000000001100100110001011101011", b"00000000000000000000000000000000"),
	(b"00000000001011101100011110110110", b"10000000000000111001101100110101"), -- -4.62726e-39 + 4.29608e-39 = -3.31184e-40
	(b"00000000001100111110000001011001", b"00000000000000000000000000000000"),
	(b"10000000001111011000101110101010", b"10000000000010011010101101010001"), -- 4.76409e-39 + -5.65207e-39 = -8.87976e-40
	(b"10000000001000100010000110110000", b"00000000000000000000000000000000"),
	(b"10000000001010011001011010000001", b"10000000010010111011100000110001"), -- -3.13449e-39 + -3.81925e-39 = -6.95374e-39
	(b"00000000011101101100010101101111", b"00000000000000000000000000000000"),
	(b"00000000001100100010000011010111", b"00000000101010001110011001000110"), -- 1.09074e-38 + 4.60356e-39 = 1.5511e-38
	(b"10000000001000011111101011110011", b"00000000000000000000000000000000"),
	(b"00000000010011100000000011100001", b"00000000001011000000010111101110"), -- -3.12059e-39 + 7.16348e-39 = 4.04289e-39
	(b"00000000000010011111111111010101", b"00000000000000000000000000000000"),
	(b"00000000000010001001011001001110", b"00000000000100101001011000100011"), -- 9.18295e-40 + 7.88603e-40 = 1.7069e-39
	(b"00000000011111001001110110100101", b"00000000000000000000000000000000"),
	(b"10000000010100110101100101001011", b"00000000001010010100010001011010"), -- 1.14442e-38 + -7.65438e-39 = 3.78978e-39
	(b"00000000010101010010000010010000", b"00000000000000000000000000000000"),
	(b"10000000001011100101000010010000", b"00000000001001101101000000000000"), -- 7.8177e-39 + -4.25333e-39 = 3.56437e-39
	(b"10000000011100011110100111100010", b"00000000000000000000000000000000"),
	(b"00000000010110111001101001011011", b"10000000000101100100111110000111"), -- -1.04613e-38 + 8.4124e-39 = -2.04891e-39
	(b"00000000010101101010001010100000", b"00000000000000000000000000000000"),
	(b"10000000010011011001100110001101", b"00000000000010010000100100010011"), -- 7.95619e-39 + -7.12642e-39 = 8.29775e-40
	(b"00000000011011111000100100111011", b"00000000000000000000000000000000"),
	(b"00000000010111101001011111001101", b"00000000110011100010000100001000"), -- 1.0243e-38 + 8.68699e-39 = 1.893e-38
	(b"00000000000010100100001010011000", b"00000000000000000000000000000000"),
	(b"10000000001000101011000110001111", b"10000000000110000110111011110111"), -- 9.42244e-40 + -3.1861e-39 = -2.24386e-39
	(b"10000000010110010010011001111111", b"00000000000000000000000000000000"),
	(b"10000000010100001111100101100010", b"10000000101010100001111111100001"), -- -8.18717e-39 + -7.4363e-39 = -1.56235e-38
	(b"00000000011111010001100110101110", b"00000000000000000000000000000000"),
	(b"00000000001001010000011000101110", b"00000000101000100001111111011100"), -- 1.14886e-38 + 3.40013e-39 = 1.48888e-38
	(b"10000000000111000110100001010110", b"00000000000000000000000000000000"),
	(b"10000000010110110001100111110001", b"10000000011101111000001001000111"), -- -2.60882e-39 + -8.36634e-39 = -1.09752e-38
	(b"00000000001111001010011100110110", b"00000000000000000000000000000000"),
	(b"10000000001010101001011001100010", b"00000000000100100001000011010100"), -- 5.57011e-39 + -3.91104e-39 = 1.65908e-39
	(b"10000000011100011110011101001011", b"00000000000000000000000000000000"),
	(b"00000000001001111000111110101110", b"10000000010010100101011110011101"), -- -1.04604e-38 + 3.63313e-39 = -6.82726e-39
	(b"00000000010100100011110000011000", b"00000000000000000000000000000000"),
	(b"10000000011101000001001100101111", b"10000000001000011101011100010111"), -- 7.55207e-39 + -1.06598e-38 = -3.10773e-39
	(b"10000000011000001000010110111100", b"00000000000000000000000000000000"),
	(b"10000000000101100100111011111010", b"10000000011101101101010010110110"), -- -8.86418e-39 + -2.04871e-39 = -1.09129e-38
	(b"10000000000000110101000111001101", b"00000000000000000000000000000000"),
	(b"00000000000100000101110011101011", b"00000000000011010000101100011110"), -- -3.04851e-40 + 1.5027e-39 = 1.19785e-39
	(b"10000000011100001111000111000111", b"00000000000000000000000000000000"),
	(b"00000000011011110110010101101110", b"10000000000000011000110001011001"), -- -1.03723e-38 + 1.02301e-38 = -1.42183e-40
	(b"00000000000001111110100110110101", b"00000000000000000000000000000000"),
	(b"10000000000101001001011001000101", b"10000000000011001010110010010000"), -- 7.26687e-40 + -1.89062e-39 = -1.16393e-39
	(b"00000000000000001010011101100101", b"00000000000000000000000000000000"),
	(b"00000000001101100110011001001111", b"00000000001101110000110110110100"), -- 6.00498e-41 + 4.99582e-39 = 5.05587e-39
	(b"10000000010101001101011011111100", b"00000000000000000000000000000000"),
	(b"00000000010111001000000001000110", b"00000000000001111010100101001010"), -- -7.7913e-39 + 8.49488e-39 = 7.03578e-40
	(b"10000000011000001000000111011100", b"00000000000000000000000000000000"),
	(b"10000000011000001000101010000001", b"10000000110000010000110001011101"), -- -8.86279e-39 + -8.86589e-39 = -1.77287e-38
	(b"00000000011010101001001101010001", b"00000000000000000000000000000000"),
	(b"00000000010011011000101100111101", b"00000000101110000001111010001110"), -- 9.78741e-39 + 7.12128e-39 = 1.69087e-38
	(b"00000000000001100100000011110000", b"00000000000000000000000000000000"),
	(b"10000000000101010101000101110110", b"10000000000011110001000010000110"), -- 5.74308e-40 + -1.95777e-39 = -1.38346e-39
	(b"10000000011110001011110110111011", b"00000000000000000000000000000000"),
	(b"10000000001011011111011001101110", b"10000000101001101011010000101001"), -- -1.10883e-38 + -4.221e-39 = -1.53093e-38
	(b"00000000010001010011110011111110", b"00000000000000000000000000000000"),
	(b"10000000010001000011001110101100", b"00000000000000010000100101010010"), -- 6.35853e-39 + -6.26335e-39 = 9.5179e-41
	(b"10000000010011101010100001010010", b"00000000000000000000000000000000"),
	(b"00000000010010001110110101000000", b"10000000000001011011101100010010"), -- -7.22355e-39 + 6.69726e-39 = -5.26286e-40
	(b"10000000011010010010110001101001", b"00000000000000000000000000000000"),
	(b"00000000010111011001010100010101", b"10000000000010111001011101010100"), -- -9.65866e-39 + 8.59418e-39 = -1.06448e-39
	(b"00000000011111110011101000100111", b"00000000000000000000000000000000"),
	(b"00000000011101100110111010100011", b"00000000111101011010100011001010"), -- 1.1684e-38 + 1.08763e-38 = 2.25602e-38
	(b"00000000000110100001101101111110", b"00000000000000000000000000000000"),
	(b"10000000000100111010100110000011", b"00000000000001100111000111111011"), -- 2.39759e-39 + -1.80568e-39 = 5.91901e-40
	(b"00000000011011011100000001011110", b"00000000000000000000000000000000"),
	(b"00000000000101001110011001000110", b"00000000100000101010011010100100"), -- 1.00791e-38 + 1.91932e-39 = 1.19984e-38
	(b"00000000001100000101111010011000", b"00000000000000000000000000000000"),
	(b"10000000000111110001011010100001", b"00000000000100010100011111110111"), -- 4.44204e-39 + -2.85502e-39 = 1.58702e-39
	(b"10000000010110111111111101101111", b"00000000000000000000000000000000"),
	(b"10000000010011001111010010110100", b"10000000101010001111010000100011"), -- -8.44866e-39 + -7.06728e-39 = -1.55159e-38
	(b"10000000000111011101111001000100", b"00000000000000000000000000000000"),
	(b"00000000001001110110110110100000", b"00000000000010011000111101011100"), -- -2.74296e-39 + 3.62091e-39 = 8.77947e-40
	(b"10000000011111001000001010010001", b"00000000000000000000000000000000"),
	(b"00000000010011010100001011111001", b"10000000001011110011111110011000"), -- -1.14344e-38 + 7.09536e-39 = -4.33908e-39
	(b"10000000000100100111101010001000", b"00000000000000000000000000000000"),
	(b"10000000010101111100011000100000", b"10000000011010100100000010101000"), -- -1.69699e-39 + -8.06076e-39 = -9.75776e-39
	(b"00000000000101101111010001111111", b"00000000000000000000000000000000"),
	(b"10000000001100011001111110000010", b"10000000000110101010101100000011"), -- 2.10809e-39 + -4.55716e-39 = -2.44907e-39
	(b"00000000011111100010000001111000", b"00000000000000000000000000000000"),
	(b"10000000001110111011100111101110", b"00000000010000100110011010001010"), -- 1.15829e-38 + -5.48499e-39 = 6.09793e-39
	(b"10000000011011001100010111000111", b"00000000000000000000000000000000"),
	(b"00000000000000001110010100111111", b"10000000011010111110000010001000"), -- -9.98918e-39 + 8.2238e-41 = -9.90694e-39
	(b"10000000010010011000001100000010", b"00000000000000000000000000000000"),
	(b"00000000000010000101011011100000", b"10000000010000010010110000100010"), -- -6.75099e-39 + 7.65849e-40 = -5.98514e-39
	(b"00000000010000001100001000101000", b"00000000000000000000000000000000"),
	(b"10000000010100101110010011111000", b"10000000000100100010001011010000"), -- 5.94712e-39 + -7.61265e-39 = -1.66553e-39
	(b"10000000011001010000111111110100", b"00000000000000000000000000000000"),
	(b"00000000000111011000111001100000", b"10000000010001111000000110010100"), -- -9.28111e-39 + 2.7143e-39 = -6.5668e-39
	(b"10000000010000111110010010111101", b"00000000000000000000000000000000"),
	(b"10000000010001100010111110001001", b"10000000100010100001010001000110"), -- -6.23503e-39 + -6.44554e-39 = -1.26806e-38
	(b"10000000001000100000110101110010", b"00000000000000000000000000000000"),
	(b"00000000011010001011001110011001", b"00000000010001101010011000100111"), -- -3.12723e-39 + 9.61532e-39 = 6.48809e-39
	(b"10000000011011101100101000001101", b"00000000000000000000000000000000"),
	(b"00000000000111011100001101111111", b"10000000010100010000011010001110"), -- -1.01744e-38 + 2.73336e-39 = -7.44103e-39
	(b"00000000001110011101101000000010", b"00000000000000000000000000000000"),
	(b"00000000010110011110110101110111", b"00000000100100111100011101111001"), -- 5.31283e-39 + 8.25855e-39 = 1.35714e-38
	(b"10000000011100011110011001010100", b"00000000000000000000000000000000"),
	(b"10000000010110000101100101101011", b"10000000110010100011111110111111"), -- -1.046e-38 + -8.1136e-39 = -1.85736e-38
	(b"00000000000101100101100111101100", b"00000000000000000000000000000000"),
	(b"10000000000110110100111010000001", b"10000000000001001111010010010101"), -- 2.05264e-39 + -2.50772e-39 = -4.55081e-40
	(b"00000000000110101000101011100011", b"00000000000000000000000000000000"),
	(b"10000000001111111111100101011010", b"10000000001001010110111001110111"), -- 2.43755e-39 + -5.87509e-39 = -3.43754e-39
	(b"00000000001010110011110101101110", b"00000000000000000000000000000000"),
	(b"10000000001010110001001101010011", b"00000000000000000010101000011011"), -- 3.97096e-39 + -3.95586e-39 = 1.51046e-41
	(b"10000000010001101000001010110011", b"00000000000000000000000000000000"),
	(b"00000000000100101010010001110010", b"10000000001100111101111001000001"), -- -6.47537e-39 + 1.71203e-39 = -4.76334e-39
	(b"00000000000011100010001001010010", b"00000000000000000000000000000000"),
	(b"00000000001110101100010101111101", b"00000000010010001110011111001111"), -- 1.29801e-39 + 5.3973e-39 = 6.69531e-39
	(b"00000000001011011001101000000110", b"00000000000000000000000000000000"),
	(b"10000000001000001001101111010110", b"00000000000011001111111000110000"), -- 4.18785e-39 + -2.99464e-39 = 1.19321e-39
	(b"00000000001001110100100000100001", b"00000000000000000000000000000000"),
	(b"10000000000100001000001001011011", b"00000000000101101100010111000110"), -- 3.60746e-39 + -1.51613e-39 = 2.09133e-39
	(b"10000000011011110111011111010101", b"00000000000000000000000000000000"),
	(b"00000000010101000001110011100011", b"10000000000110110101101011110010"), -- -1.02367e-38 + 7.72454e-39 = -2.51218e-39
	(b"10000000001010111100100001000001", b"00000000000000000000000000000000"),
	(b"10000000000010100000011010101110", b"10000000001101011100111011101111"), -- -4.02076e-39 + -9.20751e-40 = -4.94152e-39
	(b"10000000000100010001111110011000", b"00000000000000000000000000000000"),
	(b"10000000011011000011101001111111", b"10000000011111010101101000010111"), -- -1.57254e-39 + -9.93922e-39 = -1.15118e-38
	(b"10000000000000010010110100011000", b"00000000000000000000000000000000"),
	(b"00000000001100110010010001000100", b"00000000001100011111011100101100"), -- -1.08012e-40 + 4.69662e-39 = 4.58861e-39
	(b"00000000011101101100100011100010", b"00000000000000000000000000000000"),
	(b"10000000000100001110011000000010", b"00000000011001011110001011100000"), -- 1.09087e-38 + -1.55188e-39 = 9.35677e-39
	(b"00000000011110010001011101010000", b"00000000000000000000000000000000"),
	(b"00000000001000100111100010001101", b"00000000100110111000111111011101"), -- 1.11205e-38 + 3.16565e-39 = 1.42861e-38
	(b"00000000001000010100111100101100", b"00000000000000000000000000000000"),
	(b"00000000011101010000011000000010", b"00000000100101100101010100101110"), -- 3.05897e-39 + 1.07469e-38 = 1.38059e-38
	(b"10000000011001000011101110011110", b"00000000000000000000000000000000"),
	(b"10000000001100011110100011010110", b"10000000100101100010010001110100"), -- -9.20494e-39 + -4.58347e-39 = -1.37884e-38
	(b"00000000011100010011111110000101", b"00000000000000000000000000000000"),
	(b"00000000001011010110001010010110", b"00000000100111101010001000011011"), -- 1.04002e-38 + 4.16796e-39 = 1.45682e-38
	(b"00000000011100101111101010100101", b"00000000000000000000000000000000"),
	(b"00000000010000110110011010000110", b"00000000101101100110000100101011"), -- 1.05592e-38 + 6.18976e-39 = 1.67489e-38
	(b"00000000001010101101111111000010", b"00000000000000000000000000000000"),
	(b"10000000010010000111101101110101", b"10000000000111011001101110110011"), -- 3.93736e-39 + -6.65644e-39 = -2.71908e-39
	(b"10000000001001111010001001110110", b"00000000000000000000000000000000"),
	(b"00000000001101001010011010011010", b"00000000000011010000010000100100"), -- -3.63986e-39 + 4.83521e-39 = 1.19535e-39
	(b"00000000011110111101010011100100", b"00000000000000000000000000000000"),
	(b"10000000001000001110100011001001", b"00000000010110101110110000011011"), -- 1.13721e-38 + -3.02224e-39 = 8.34989e-39
	(b"10000000010101011111111110110110", b"00000000000000000000000000000000"),
	(b"10000000011111001010111001111101", b"10000000110100101010111000110011"), -- -7.89775e-39 + -1.14502e-38 = -1.93479e-38
	(b"10000000011010000110100000010001", b"00000000000000000000000000000000"),
	(b"10000000011101010110010101110000", b"10000000110111011100110110000001"), -- -9.58822e-39 + -1.07811e-38 = -2.03694e-38
	(b"10000000000000111010000111100110", b"00000000000000000000000000000000"),
	(b"00000000000011011111011000101001", b"00000000000010100101010001000011"), -- -3.33585e-40 + 1.28217e-39 = 9.48582e-40
	(b"10000000000100100011000100000101", b"00000000000000000000000000000000"),
	(b"10000000011001000000000100110110", b"10000000011101100011001000111011"), -- -1.67062e-39 + -9.18398e-39 = -1.08546e-38
	(b"00000000011101100101010011011011", b"00000000000000000000000000000000"),
	(b"10000000000001111100111011100011", b"00000000011011101000010111111000"), -- 1.0867e-38 + -7.17065e-40 = 1.015e-38
	(b"10000000010111110111010110101000", b"00000000000000000000000000000000"),
	(b"00000000011010010000111110010010", b"00000000000010011001100111101010"), -- -8.76658e-39 + 9.64831e-39 = 8.81733e-40
	(b"10000000011110011101110101111001", b"00000000000000000000000000000000"),
	(b"10000000011000001100011111110001", b"10000000110110101010010101101010"), -- -1.11915e-38 + -8.88793e-39 = -2.00795e-38
	(b"10000000001100111101011110010111", b"00000000000000000000000000000000"),
	(b"00000000010011101011010111101000", b"00000000000110101101111001010001"), -- -4.76095e-39 + 7.22842e-39 = 2.46747e-39
	(b"00000000010000011111111001111101", b"00000000000000000000000000000000"),
	(b"10000000000111101001110110110010", b"00000000001000110110000011001011"), -- 6.0606e-39 + -2.81164e-39 = 3.24897e-39
	(b"10000000000011011001010100101111", b"00000000000000000000000000000000"),
	(b"10000000010110001010100000000000", b"10000000011001100011110100101111"), -- -1.24738e-39 + -8.14179e-39 = -9.38917e-39
	(b"10000000010110001100110111011101", b"00000000000000000000000000000000"),
	(b"10000000010101100100000110001110", b"10000000101011110000111101101011"), -- -8.15537e-39 + -7.92137e-39 = -1.60767e-38
	(b"10000000010101110101101001011011", b"00000000000000000000000000000000"),
	(b"00000000000001000001001001100100", b"10000000010100110100011111110111"), -- -8.0221e-39 + 3.73939e-40 = -7.64816e-39
	(b"00000000000011011010110101100011", b"00000000000000000000000000000000"),
	(b"10000000010110100010101001000000", b"10000000010011000111110011011101"), -- 1.25606e-39 + -8.28035e-39 = -7.02429e-39
	(b"10000000000010011001110111010011", b"00000000000000000000000000000000"),
	(b"10000000010000111110011110000011", b"10000000010011011000010101010110"), -- -8.83136e-40 + -6.23603e-39 = -7.11917e-39
	(b"10000000011111001001100111010010", b"00000000000000000000000000000000"),
	(b"00000000011000001010001100010011", b"10000000000110111111011010111111"), -- -1.14428e-38 + 8.87471e-39 = -2.56807e-39
	(b"00000000001100000001110011101101", b"00000000000000000000000000000000"),
	(b"10000000011101111001010000000110", b"10000000010001110111011100011001"), -- 4.41848e-39 + -1.09815e-38 = -6.56304e-39
	(b"00000000000011111111101101001101", b"00000000000000000000000000000000"),
	(b"00000000000100010000101101011111", b"00000000001000010000011010101100"), -- 1.46768e-39 + 1.56528e-39 = 3.03296e-39
	(b"10000000001000010101110000010000", b"00000000000000000000000000000000"),
	(b"10000000010011000010110110010000", b"10000000011011011000100110100000"), -- -3.0636e-39 + -6.99584e-39 = -1.00594e-38
	(b"10000000000010000100110111111101", b"00000000000000000000000000000000"),
	(b"10000000011011011010110000110000", b"10000000011101011111101000101101"), -- -7.62661e-40 + -1.00718e-38 = -1.08345e-38
	(b"10000000010110011100101000110110", b"00000000000000000000000000000000"),
	(b"10000000001010100111010110101110", b"10000000100001000011111111100100"), -- -8.2459e-39 + -3.89931e-39 = -1.21452e-38
	(b"10000000001110111110001000011011", b"00000000000000000000000000000000"),
	(b"10000000011001011000110001011100", b"10000000101000010110111001110111"), -- -5.49941e-39 + -9.32574e-39 = -1.48251e-38
	(b"10000000010110101111110100101110", b"00000000000000000000000000000000"),
	(b"00000000000001100011001000100010", b"10000000010101001100101100001100"), -- -8.35602e-39 + 5.68997e-40 = -7.78702e-39
	(b"00000000001001111110000001100110", b"00000000000000000000000000000000"),
	(b"10000000011000000011110111111001", b"10000000001110000101110110010011"), -- 3.66208e-39 + -8.83844e-39 = -5.17636e-39
	(b"10000000000010001101101111110001", b"00000000000000000000000000000000"),
	(b"00000000000011001010010100110000", b"00000000000000111100100100111111"), -- -8.13584e-40 + 1.16128e-39 = 3.477e-40
	(b"10000000000110011101111100011000", b"00000000000000000000000000000000"),
	(b"10000000010010101011111000001011", b"10000000011001001001110100100011"), -- -2.37592e-39 + -6.864e-39 = -9.23992e-39
	(b"10000000000010101100110010010010", b"00000000000000000000000000000000"),
	(b"10000000011000011101010100110111", b"10000000011011001010000111001001"), -- -9.91741e-40 + -8.98453e-39 = -9.97627e-39
	(b"00000000011001010111100101101011", b"00000000000000000000000000000000"),
	(b"10000000000110100000000001101000", b"00000000010010110111100100000011"), -- 9.31894e-39 + -2.38787e-39 = 6.93107e-39
	(b"10000000000010110110110110011101", b"00000000000000000000000000000000"),
	(b"10000000000011001100110111110001", b"10000000000110000011101110001110"), -- -1.04951e-39 + -1.1759e-39 = -2.22542e-39
	(b"10000000000010110010110101111101", b"00000000000000000000000000000000"),
	(b"10000000011010011000110001000000", b"10000000011101001011100110111101"), -- -1.02651e-39 + -9.69304e-39 = -1.07195e-38
	(b"00000000011011111000101011111001", b"00000000000000000000000000000000"),
	(b"00000000011110010000010010000000", b"00000000111010001000111101111001"), -- 1.02436e-38 + 1.11137e-38 = 2.13573e-38
	(b"00000000011100000000111001101010", b"00000000000000000000000000000000"),
	(b"10000000000011111001001110100100", b"00000000011000000111101011000110"), -- 1.02907e-38 + -1.4305e-39 = 8.86025e-39
	(b"00000000001111011000001010101011", b"00000000000000000000000000000000"),
	(b"10000000010000000000011010010011", b"10000000000000101000001111101000"), -- 5.64884e-39 + -5.87983e-39 = -2.3099e-40
	(b"10000000000000000101001111011010", b"00000000000000000000000000000000"),
	(b"10000000010011101111011100111000", b"10000000010011110100101100010010"), -- -3.00803e-41 + -7.25185e-39 = -7.28193e-39
	(b"10000000010001011001011101101101", b"00000000000000000000000000000000"),
	(b"00000000011000001010101100111110", b"00000000000110110001001111010001"), -- -6.39097e-39 + 8.87764e-39 = 2.48667e-39
	(b"10000000011100011100001110100001", b"00000000000000000000000000000000"),
	(b"00000000010101010000011111011101", b"10000000000111001011101111000100"), -- -1.04476e-38 + 7.80884e-39 = -2.63875e-39
	(b"00000000011110010011110010010011", b"00000000000000000000000000000000"),
	(b"10000000010101000010010110010000", b"00000000001001010001011100000011"), -- 1.11338e-38 + -7.72766e-39 = 3.40617e-39
	(b"10000000000001011010100001111101", b"00000000000000000000000000000000"),
	(b"00000000010000110000100111001011", b"00000000001111010110000101001110"), -- -5.1962e-40 + 6.15649e-39 = 5.63687e-39
	(b"10000000010110000010000000000000", b"00000000000000000000000000000000"),
	(b"00000000011110100001111000111111", b"00000000001000011111111000111111"), -- -8.093e-39 + 1.12148e-38 = 3.12178e-39
	(b"10000000011111101011101101011111", b"00000000000000000000000000000000"),
	(b"00000000001110100101010101111101", b"10000000010001000110010111100010"), -- -1.16385e-38 + 5.35713e-39 = -6.28136e-39
	(b"10000000001101111110001110110011", b"00000000000000000000000000000000"),
	(b"10000000010010111110111001011011", b"10000000100000111101001000001110"), -- -5.13264e-39 + -6.97317e-39 = -1.21058e-38
	(b"10000000001010110110011101101011", b"00000000000000000000000000000000"),
	(b"10000000011100101001111101110100", b"10000000100111100000011011011111"), -- -3.98603e-39 + -1.05264e-38 = -1.45125e-38
	(b"00000000011000110010111101111100", b"00000000000000000000000000000000"),
	(b"00000000000110110110101010100000", b"00000000011111101001101000011100"), -- 9.10875e-39 + 2.51781e-39 = 1.16266e-38
	(b"10000000011001000100110111110100", b"00000000000000000000000000000000"),
	(b"10000000011001100110101011110111", b"10000000110010101011100011101011"), -- -9.21151e-39 + -9.40559e-39 = -1.86171e-38
	(b"00000000011101010001011001100111", b"00000000000000000000000000000000"),
	(b"10000000000110000001100001000010", b"00000000010111001111111000100101"), -- 1.07528e-38 + -2.21275e-39 = 8.54004e-39
	(b"00000000000000111110010001100111", b"00000000000000000000000000000000"),
	(b"00000000000001101101110100110011", b"00000000000010101100000110011010"), -- 3.57442e-40 + 6.30364e-40 = 9.87806e-40
	(b"10000000001110111111010010011101", b"00000000000000000000000000000000"),
	(b"00000000011001010100100001111111", b"00000000001010010101001111100010"), -- -5.50604e-39 + 9.30139e-39 = 3.79535e-39
	(b"10000000010101000101001101101011", b"00000000000000000000000000000000"),
	(b"00000000010000000111010001000100", b"10000000000100111101111100100111"), -- -7.74411e-39 + 5.91918e-39 = -1.82493e-39
	(b"00000000010100110001100111101001", b"00000000000000000000000000000000"),
	(b"00000000011101101101100000100101", b"00000000110010011111001000001110"), -- 7.63164e-39 + 1.09141e-38 = 1.85458e-38
	(b"00000000010001100010101110101011", b"00000000000000000000000000000000"),
	(b"00000000000001110100010010000001", b"00000000010011010111000000101100"), -- 6.44415e-39 + 6.67423e-40 = 7.11157e-39
	(b"00000000001101100100011001101010", b"00000000000000000000000000000000"),
	(b"10000000010010100101000100101110", b"10000000000101000000101011000100"), -- 4.98438e-39 + -6.82495e-39 = -1.84057e-39
	(b"00000000001000011110011110010100", b"00000000000000000000000000000000"),
	(b"00000000010110011010010111010110", b"00000000011110111000110101101010"), -- 3.11365e-39 + 8.23285e-39 = 1.13465e-38
	(b"00000000010111111001010111101000", b"00000000000000000000000000000000"),
	(b"00000000000101100101111101111011", b"00000000011101011111010101100011"), -- 8.77815e-39 + 2.05463e-39 = 1.08328e-38
	(b"00000000011010101110111111110001", b"00000000000000000000000000000000"),
	(b"00000000010100011110010011001000", b"00000000101111001101010010111001"), -- 9.82064e-39 + 7.52075e-39 = 1.73414e-38
	(b"00000000011100010001011010000011", b"00000000000000000000000000000000"),
	(b"00000000001100110010110000011100", b"00000000101001000100001010011111"), -- 1.03855e-38 + 4.69943e-39 = 1.50849e-38
	(b"10000000010111111100110110001000", b"00000000000000000000000000000000"),
	(b"00000000000000010110011111000100", b"10000000010111100110010111000100"), -- -8.7981e-39 + 1.2906e-40 = -8.66904e-39
	(b"00000000001111001011111100101110", b"00000000000000000000000000000000"),
	(b"10000000000100101101111001011011", b"00000000001010011110000011010011"), -- 5.57871e-39 + -1.73281e-39 = 3.84591e-39
	(b"00000000010000010000001101100000", b"00000000000000000000000000000000"),
	(b"00000000000100101101101110000101", b"00000000010100111101111011100101"), -- 5.97052e-39 + 1.73179e-39 = 7.70231e-39
	(b"10000000011100100001100001110111", b"00000000000000000000000000000000"),
	(b"00000000001111100010100100111000", b"10000000001100111110111100111111"), -- -1.0478e-38 + 5.70859e-39 = -4.76944e-39
	(b"00000000010100100010010000001010", b"00000000000000000000000000000000"),
	(b"00000000000011001101010010100110", b"00000000010111101111100010110000"), -- 7.54344e-39 + 1.17831e-39 = 8.72175e-39
	(b"00000000000110010001000010010000", b"00000000000000000000000000000000"),
	(b"10000000011100001000011100001010", b"10000000010101110111011001111010"), -- 2.30183e-39 + -1.0334e-38 = -8.03219e-39
	(b"10000000010101010100110100110110", b"00000000000000000000000000000000"),
	(b"00000000001000011101000100111001", b"10000000001100110111101111111101"), -- -7.83372e-39 + 3.10563e-39 = -4.72809e-39
	(b"10000000010001101100001101101111", b"00000000000000000000000000000000"),
	(b"10000000001100100011111101111101", b"10000000011110010000001011101100"), -- -6.49859e-39 + -4.61455e-39 = -1.11131e-38
	(b"00000000001000000010101011111100", b"00000000000000000000000000000000"),
	(b"10000000011101101100111011101000", b"10000000010101101010001111101100"), -- 2.95416e-39 + -1.09108e-38 = -7.95666e-39
	(b"00000000001011001100001000100110", b"00000000000000000000000000000000"),
	(b"10000000000011001011100000111101", b"00000000001000000000100111101001"), -- 4.11041e-39 + -1.16812e-39 = 2.94229e-39
	(b"00000000010000001001011001110000", b"00000000000000000000000000000000"),
	(b"10000000000001100110010101110011", b"00000000001110100011000011111101"), -- 5.93144e-39 + -5.87406e-40 = 5.34403e-39
	(b"00000000001110010110001000010111", b"00000000000000000000000000000000"),
	(b"00000000010111000000000010110001", b"00000000100101010110001011001000"), -- 5.26981e-39 + 8.44911e-39 = 1.37189e-38
	(b"10000000000110011100111100110000", b"00000000000000000000000000000000"),
	(b"00000000010011001001111010110011", b"00000000001100101100111110000011"), -- -2.37021e-39 + 7.03643e-39 = 4.66622e-39
	(b"00000000011110000110111111011000", b"00000000000000000000000000000000"),
	(b"00000000010110011010110100101001", b"00000000110100100001110100000001"), -- 1.10604e-38 + 8.23548e-39 = 1.92959e-38
	(b"00000000000001010001111100100110", b"00000000000000000000000000000000"),
	(b"10000000001010001011010111001000", b"10000000001000111001011010100010"), -- 4.70351e-40 + -3.73863e-39 = -3.26828e-39
	(b"10000000011110000001001101111010", b"00000000000000000000000000000000"),
	(b"10000000001000110001001000011001", b"10000000100110110010010110010011"), -- -1.10272e-38 + -3.22073e-39 = -1.4248e-38
	(b"00000000000100011010100110001000", b"00000000000000000000000000000000"),
	(b"00000000001101101000010001011110", b"00000000010010000010110111100110"), -- 1.62202e-39 + 5.0066e-39 = 6.62862e-39
	(b"00000000001101111101110011111011", b"00000000000000000000000000000000"),
	(b"00000000001001010100101111110110", b"00000000010111010010100011110001"), -- 5.13023e-39 + 3.42516e-39 = 8.55539e-39
	(b"00000000011101000001111010011000", b"00000000000000000000000000000000"),
	(b"10000000010000011010011111010110", b"00000000001100100111011011000010"), -- 1.06639e-38 + -6.02952e-39 = 4.63438e-39
	(b"10000000000100011100111101101001", b"00000000000000000000000000000000"),
	(b"00000000010101101111111101010001", b"00000000010001010010111111101000"), -- -1.63561e-39 + 7.98944e-39 = 6.35383e-39
	(b"00000000001000100100010110111001", b"00000000000000000000000000000000"),
	(b"10000000010010111100010111011011", b"10000000001010011000000000100010"), -- 3.14742e-39 + -6.95864e-39 = -3.81122e-39
	(b"00000000010010010101000001101000", b"00000000000000000000000000000000"),
	(b"10000000001001000011101111110001", b"00000000001001010001010001110111"), -- 6.73284e-39 + -3.32758e-39 = 3.40525e-39
	(b"10000000011011001010111111010011", b"00000000000000000000000000000000"),
	(b"00000000001000111110001000100001", b"10000000010010001100110110110010"), -- -9.98131e-39 + 3.29536e-39 = -6.68595e-39
	(b"00000000000011010101110001010000", b"00000000000000000000000000000000"),
	(b"10000000010110101110101000000000", b"10000000010011011000110110110000"), -- 1.22698e-39 + -8.34914e-39 = -7.12216e-39
	(b"10000000001001111001100111100011", b"00000000000000000000000000000000"),
	(b"10000000000101010010001011101101", b"10000000001111001011110011010000"), -- -3.63679e-39 + -1.94107e-39 = -5.57786e-39
	(b"00000000000101101110010110101001", b"00000000000000000000000000000000"),
	(b"10000000000001011100101111010100", b"00000000000100010001100111010101"), -- 2.10277e-39 + -5.32297e-40 = 1.57047e-39
	(b"00000000010110100111000001000110", b"00000000000000000000000000000000"),
	(b"00000000011111000011001110110000", b"00000000110101101010001111110110"), -- 8.30547e-39 + 1.14061e-38 = 1.97116e-38
	(b"10000000001110011000110001011001", b"00000000000000000000000000000000"),
	(b"10000000000110111101001001001101", b"10000000010101010101111010100110"), -- -5.28497e-39 + -2.555e-39 = -7.83997e-39
	(b"10000000000111001001011100001000", b"00000000000000000000000000000000"),
	(b"10000000000110011101101101001011", b"10000000001101100111001001010011"), -- -2.62557e-39 + -2.37455e-39 = -5.00013e-39
	(b"10000000011111000101010101110110", b"00000000000000000000000000000000"),
	(b"00000000010000000111011101100001", b"10000000001110111101111000010101"), -- -1.14183e-38 + 5.9203e-39 = -5.49796e-39
	(b"10000000011110100100100000110011", b"00000000000000000000000000000000"),
	(b"10000000010101110110100010100011", b"10000000110100011011000011010110"), -- -1.12298e-38 + -8.02722e-39 = -1.92571e-38
	(b"00000000011111101101000100011100", b"00000000000000000000000000000000"),
	(b"00000000010110010001110111000101", b"00000000110101111110111011100001"), -- 1.16463e-38 + 8.18404e-39 = 1.98303e-38
	(b"00000000000000100011011010011101", b"00000000000000000000000000000000"),
	(b"10000000001110001011001100000010", b"10000000001101100111110001100101"), -- 2.03263e-40 + -5.207e-39 = -5.00374e-39
	(b"10000000010010111110000111110111", b"00000000000000000000000000000000"),
	(b"10000000010110010001011001001111", b"10000000101001001111100001000110"), -- -6.96872e-39 + -8.18136e-39 = -1.51501e-38
	(b"00000000000011110001110101010101", b"00000000000000000000000000000000"),
	(b"10000000011001011001100010110000", b"10000000010101100111101101011011"), -- 1.38805e-39 + -9.33016e-39 = -7.9421e-39
	(b"00000000011101100011101010101001", b"00000000000000000000000000000000"),
	(b"00000000010011110110001001100010", b"00000000110001011001110100001011"), -- 1.08576e-38 + 7.2903e-39 = 1.81479e-38
	(b"00000000011000010110111100100110", b"00000000000000000000000000000000"),
	(b"10000000000011010011000111110011", b"00000000010101000011110100110011"), -- 8.94792e-39 + -1.21178e-39 = 7.73614e-39
	(b"00000000000111100000001111010100", b"00000000000000000000000000000000"),
	(b"10000000000111110010110010001110", b"10000000000000010010100010111010"), -- 2.75644e-39 + -2.86288e-39 = -1.06445e-40
	(b"00000000010111001110011101000101", b"00000000000000000000000000000000"),
	(b"00000000001011110010001100001100", b"00000000100011000000101001010001"), -- 8.53183e-39 + 4.32884e-39 = 1.28607e-38
	(b"00000000001101111111101111100010", b"00000000000000000000000000000000"),
	(b"00000000011010000100011011010100", b"00000000101000000100001010110110"), -- 5.14131e-39 + 9.5763e-39 = 1.47176e-38
	(b"10000000010111100111110100100111", b"00000000000000000000000000000000"),
	(b"10000000001011101000001010010101", b"10000000100011001111111110111100"), -- -8.67743e-39 + -4.27128e-39 = -1.29487e-38
	(b"00000000010011100010001110001111", b"00000000000000000000000000000000"),
	(b"00000000001010001001000010100110", b"00000000011101101011010000110101"), -- 7.17592e-39 + 3.72531e-39 = 1.09012e-38
	(b"00000000011101001010110100110000", b"00000000000000000000000000000000"),
	(b"10000000011101011011001010000011", b"10000000000000010000010101010011"), -- 1.0715e-38 + -1.08088e-38 = -9.37455e-41
	(b"10000000001010110000010100010010", b"00000000000000000000000000000000"),
	(b"00000000001001101011000100100011", b"10000000000001000101001111101111"), -- -3.95075e-39 + 3.55329e-39 = -3.97452e-40
	(b"10000000011101101000001000000001", b"00000000000000000000000000000000"),
	(b"00000000000010001001011001101110", b"10000000011011011110101110010011"), -- -1.08832e-38 + 7.88648e-40 = -1.00946e-38
	(b"10000000010111010010101000001100", b"00000000000000000000000000000000"),
	(b"00000000001100001011001111100001", b"10000000001011000111011000101011"), -- -8.55578e-39 + 4.47263e-39 = -4.08315e-39
	(b"10000000001011001110001100010001", b"00000000000000000000000000000000"),
	(b"00000000010000010100101100011100", b"00000000000101000110100000001011"), -- -4.12222e-39 + 5.99625e-39 = 1.87403e-39
	(b"00000000000101111001100100110110", b"00000000000000000000000000000000"),
	(b"10000000000111011100110101000001", b"10000000000001100011010000001011"), -- 2.16718e-39 + -2.73686e-39 = -5.69682e-40
	(b"10000000010110011011011100100000", b"00000000000000000000000000000000"),
	(b"10000000010000001011000110000101", b"10000000100110100110100010100101"), -- -8.23905e-39 + -5.94115e-39 = -1.41802e-38
	(b"00000000010011001110111100010010", b"00000000000000000000000000000000"),
	(b"10000000001000010001110010110001", b"00000000001010111101001001100001"), -- 7.06526e-39 + -3.04086e-39 = 4.0244e-39
	(b"00000000011111000011101111011001", b"00000000000000000000000000000000"),
	(b"10000000001101101000111010101111", b"00000000010001011010110100101010"), -- 1.14091e-38 + -5.0103e-39 = 6.39877e-39
	(b"00000000010100000000010111011011", b"00000000000000000000000000000000"),
	(b"10000000010001010100110110011111", b"00000000000010101011100000111100"), -- 7.34894e-39 + -6.36449e-39 = 9.84446e-40
	(b"00000000000101001010101111101011", b"00000000000000000000000000000000"),
	(b"00000000010011011011111010111101", b"00000000011000100110101010101000"), -- 1.89838e-39 + 7.13976e-39 = 9.03814e-39
	(b"10000000011100010010011101111111", b"00000000000000000000000000000000"),
	(b"00000000010110101011101100000011", b"10000000000101100110110001111100"), -- -1.03916e-38 + 8.33228e-39 = -2.0593e-39
	(b"00000000000111110001001011101010", b"00000000000000000000000000000000"),
	(b"10000000011110100110011110011110", b"10000000010110110101010010110100"), -- 2.85369e-39 + -1.12411e-38 = -8.38742e-39
	(b"10000000001101001001001101001110", b"00000000000000000000000000000000"),
	(b"10000000011011000100000110001100", b"10000000101000001101010011011010"), -- -4.82829e-39 + -9.94175e-39 = -1.477e-38
	(b"00000000010011011110010111100000", b"00000000000000000000000000000000"),
	(b"10000000001111101010001111001000", b"00000000000011110100001000011000"), -- 7.1538e-39 + -5.75255e-39 = 1.40124e-39
	(b"10000000011111111100101011110111", b"00000000000000000000000000000000"),
	(b"10000000011011000001001000101111", b"10000000111010111101110100100110"), -- -1.17359e-38 + -9.92476e-39 = -2.16607e-38
	(b"10000000011101000011011010010011", b"00000000000000000000000000000000"),
	(b"10000000000101101001110110010011", b"10000000100010101101010000100110"), -- -1.06725e-38 + -2.07691e-39 = -1.27494e-38
	(b"00000000010100111000110010010010", b"00000000000000000000000000000000"),
	(b"00000000000001111011000011011000", b"00000000010110110011110101101010"), -- 7.67277e-39 + 7.06288e-40 = 8.37906e-39
	(b"10000000001010100100000000111100", b"00000000000000000000000000000000"),
	(b"00000000001101011000111111010000", b"00000000000010110100111110010100"), -- -3.88013e-39 + 4.91887e-39 = 1.03874e-39
	(b"10000000001100100110011100111111", b"00000000000000000000000000000000"),
	(b"00000000001100110011100101101100", b"00000000000000001101001000101101"), -- -4.62881e-39 + 4.70421e-39 = 7.53969e-41
	(b"10000000011101000011100111101011", b"00000000000000000000000000000000"),
	(b"10000000000010111110100110011010", b"10000000100000000010001110000101"), -- -1.06737e-38 + -1.09399e-39 = -1.17677e-38
	(b"00000000001110100110010000110011", b"00000000000000000000000000000000"),
	(b"10000000001000011101100010111111", b"00000000000110001000101101110100"), -- 5.3624e-39 + -3.10833e-39 = 2.25408e-39
	(b"00000000000001000111010101111010", b"00000000000000000000000000000000"),
	(b"00000000011111100010111000110100", b"00000000100000101010001110101110"), -- 4.09485e-40 + 1.15878e-38 = 1.19973e-38
	(b"00000000001111010100111101100111", b"00000000000000000000000000000000"),
	(b"10000000010010100110001100110100", b"10000000000011010001001111001101"), -- 5.63045e-39 + -6.83141e-39 = -1.20096e-39
	(b"10000000011000100000110010111100", b"00000000000000000000000000000000"),
	(b"00000000001110001001100100110111", b"10000000001010010111001110000101"), -- -9.00445e-39 + 5.19775e-39 = -3.8067e-39
	(b"00000000001110001000010010101110", b"00000000000000000000000000000000"),
	(b"10000000000011111011010000001000", b"00000000001010001101000010100110"), -- 5.19038e-39 + -1.44212e-39 = 3.74827e-39
	(b"10000000001001010100110010111100", b"00000000000000000000000000000000"),
	(b"00000000011111001011001001000100", b"00000000010101110110010110001000"), -- -3.42544e-39 + 1.14516e-38 = 8.02611e-39
	(b"00000000000000001011110010101111", b"00000000000000000000000000000000"),
	(b"00000000000100111000010010111001", b"00000000000101000100000101101000"), -- 6.76869e-41 + 1.79249e-39 = 1.86017e-39
	(b"00000000000110110110011001110110", b"00000000000000000000000000000000"),
	(b"10000000001111101011100110110011", b"10000000001000110101001100111101"), -- 2.51631e-39 + -5.76042e-39 = -3.2441e-39
	(b"10000000000000111101011111110101", b"00000000000000000000000000000000"),
	(b"10000000000001101101001100010000", b"10000000000010101010101100000101"), -- -3.52977e-40 + -6.26728e-40 = -9.79705e-40
	(b"10000000011110110011011011101110", b"00000000000000000000000000000000"),
	(b"10000000000001101110111010010111", b"10000000100000100010010110000101"), -- -1.13155e-38 + -6.36603e-40 = -1.19521e-38
	(b"10000000011111001110001001000000", b"00000000000000000000000000000000"),
	(b"10000000001110101101010010010001", b"10000000101101111011011011010001"), -- -1.14688e-38 + -5.40271e-39 = -1.68715e-38
	(b"10000000001010001000000110100110", b"00000000000000000000000000000000"),
	(b"00000000010000011111011111000001", b"00000000000110010111011000011011"), -- -3.71993e-39 + 6.05818e-39 = 2.33826e-39
	(b"10000000011100110110011010101101", b"00000000000000000000000000000000"),
	(b"10000000001110000110110000011011", b"10000000101010111101001011001000"), -- -1.05979e-38 + -5.18157e-39 = -1.57795e-38
	(b"10000000000101000101101011101100", b"00000000000000000000000000000000"),
	(b"00000000001110111000001011111010", b"00000000001001110010100000001110"), -- -1.86933e-39 + 5.46528e-39 = 3.59595e-39
	(b"10000000000101110000100001111110", b"00000000000000000000000000000000"),
	(b"10000000000000000111100010001110", b"10000000000101111000000100001100"), -- -2.11526e-39 + -4.32469e-41 = -2.15851e-39
	(b"10000000011000011110010011000100", b"00000000000000000000000000000000"),
	(b"00000000011001101110110001111100", b"00000000000001010000011110111000"), -- -8.99011e-39 + 9.45206e-39 = 4.61946e-40
	(b"10000000011000100000011000010100", b"00000000000000000000000000000000"),
	(b"10000000001010100100111110111010", b"10000000100011000101010111001110"), -- -9.00206e-39 + -3.88569e-39 = -1.28878e-38
	(b"00000000001101010010011100000111", b"00000000000000000000000000000000"),
	(b"10000000001111011101100000111000", b"10000000000010001011000100110001"), -- 4.88128e-39 + -5.67953e-39 = -7.98248e-40
	(b"10000000010001011110010000111010", b"00000000000000000000000000000000"),
	(b"00000000010100000110010001110111", b"00000000000010101000000000111101"), -- -6.41852e-39 + 7.38288e-39 = 9.64358e-40
	(b"10000000000101001001011000000101", b"00000000000000000000000000000000"),
	(b"00000000011101010001101111011101", b"00000000011000001000010111011000"), -- -1.89053e-39 + 1.07547e-38 = 8.86422e-39
	(b"10000000000111100100010111010010", b"00000000000000000000000000000000"),
	(b"10000000010110100101001011011110", b"10000000011110001001100010110000"), -- -2.78011e-39 + -8.29492e-39 = -1.1075e-38
	(b"10000000010110111001111001111101", b"00000000000000000000000000000000"),
	(b"10000000011000101010101010000111", b"10000000101111100100100100000100"), -- -8.41389e-39 + -9.06105e-39 = -1.74749e-38
	(b"00000000010101001000110101000011", b"00000000000000000000000000000000"),
	(b"10000000001110010011011010011110", b"00000000000110110101011010100101"), -- 7.76486e-39 + -5.25422e-39 = 2.51064e-39
	(b"10000000000110000001101101010010", b"00000000000000000000000000000000"),
	(b"10000000001110001010001101101011", b"10000000010100001011111010111101"), -- -2.21385e-39 + -5.20141e-39 = -7.41526e-39
	(b"10000000010111100001001001001001", b"00000000000000000000000000000000"),
	(b"10000000001000101000001110011011", b"10000000100000001001010111100100"), -- -8.6391e-39 + -3.16962e-39 = -1.18087e-38
	(b"00000000000100010101101111010110", b"00000000000000000000000000000000"),
	(b"00000000011101100011011000110011", b"00000000100001111001001000001001"), -- 1.59415e-39 + 1.0856e-38 = 1.24502e-38
	(b"10000000011000000101011010100000", b"00000000000000000000000000000000"),
	(b"10000000011100110011001110011101", b"10000000110100111000101000111101"), -- -8.84728e-39 + -1.05796e-38 = -1.94269e-38
	(b"00000000010000011000111000111110", b"00000000000000000000000000000000"),
	(b"10000000010011001011101101011010", b"10000000000010110010110100011100"), -- 6.02033e-39 + -7.04671e-39 = -1.02637e-39
	(b"00000000000111001101010010010101", b"00000000000000000000000000000000"),
	(b"00000000001000101100101101101001", b"00000000001111111001111111111110"), -- 2.64765e-39 + 3.19538e-39 = 5.84303e-39
	(b"10000000001011100010010110110111", b"00000000000000000000000000000000"),
	(b"10000000011010001000000010001111", b"10000000100101101010011001000110"), -- -4.23796e-39 + -9.59701e-39 = -1.3835e-38
	(b"10000000011010011111000100110000", b"00000000000000000000000000000000"),
	(b"00000000000110000100111111011100", b"10000000010100011010000101010100"), -- -9.72925e-39 + 2.2327e-39 = -7.49655e-39
	(b"00000000000111000001110011010110", b"00000000000000000000000000000000"),
	(b"10000000010100011100000101101001", b"10000000001101011010010010010011"), -- 2.58174e-39 + -7.50806e-39 = -4.92632e-39
	(b"10000000000110101001100010011110", b"00000000000000000000000000000000"),
	(b"10000000001001111101011111011011", b"10000000010000100111000001111001"), -- -2.44247e-39 + -3.65902e-39 = -6.10149e-39
	(b"00000000000011100100110111111110", b"00000000000000000000000000000000"),
	(b"00000000010111101101110101101011", b"00000000011011010010101101101001"), -- 1.31368e-39 + 8.71197e-39 = 1.00256e-38
	(b"00000000001111111000011001001111", b"00000000000000000000000000000000"),
	(b"00000000000111111111010110010111", b"00000000010111110111101111100110"), -- 5.83382e-39 + 2.935e-39 = 8.76882e-39
	(b"10000000011011011111010100110000", b"00000000000000000000000000000000"),
	(b"10000000011101100100101000101000", b"10000000111001000011111101011000"), -- -1.0098e-38 + -1.08632e-38 = -2.09612e-38
	(b"00000000010010100110110010110110", b"00000000000000000000000000000000"),
	(b"10000000011011010011111001011100", b"10000000001000101101000110100110"), -- 6.83482e-39 + -1.00324e-38 = -3.19761e-39
	(b"00000000010110000011001000001010", b"00000000000000000000000000000000"),
	(b"10000000001000110111111000111111", b"00000000001101001011001111001011"), -- 8.09947e-39 + -3.25953e-39 = 4.83994e-39
	(b"00000000011101110101111101010000", b"00000000000000000000000000000000"),
	(b"00000000001000001001110000111101", b"00000000100101111111101110001101"), -- 1.09626e-38 + 2.99478e-39 = 1.39574e-38
	(b"10000000000001111100000011100110", b"00000000000000000000000000000000"),
	(b"00000000011100000001101001101111", b"00000000011010000101100110001001"), -- -7.12047e-40 + 1.02951e-38 = 9.58301e-39
	(b"10000000011110110011011110000100", b"00000000000000000000000000000000"),
	(b"00000000000001001011001100000001", b"10000000011101101000010010000011"), -- -1.13157e-38 + 4.31556e-40 = -1.08841e-38
	(b"10000000001110111110111010010000", b"00000000000000000000000000000000"),
	(b"10000000011010001100000101001110", b"10000000101001001010111111011110"), -- -5.50387e-39 + -9.62024e-39 = -1.51241e-38
	(b"10000000011101001110000110001011", b"00000000000000000000000000000000"),
	(b"00000000011110101001111001111010", b"00000000000001011011110011101111"), -- -1.07338e-38 + 1.12608e-38 = 5.26954e-40
	(b"10000000001110011110010110000000", b"00000000000000000000000000000000"),
	(b"00000000011011000000110000010000", b"00000000001100100010011010010000"), -- -5.31695e-39 + 9.92256e-39 = 4.60561e-39
	(b"00000000000111010011000011110000", b"00000000000000000000000000000000"),
	(b"00000000011101000010011100001001", b"00000000100100010101011111111001"), -- 2.68078e-39 + 1.06669e-38 = 1.33477e-38
	(b"00000000011101110011001111010010", b"00000000000000000000000000000000"),
	(b"00000000011011101000101001110101", b"00000000111001011011111001000111"), -- 1.0947e-38 + 1.01516e-38 = 2.10986e-38
	(b"10000000010111010101000110101100", b"00000000000000000000000000000000"),
	(b"10000000000100101011011111101011", b"10000000011100000000100110010111"), -- -8.57e-39 + -1.71902e-39 = -1.0289e-38
	(b"00000000011011011100000110101101", b"00000000000000000000000000000000"),
	(b"10000000001001110101011010110011", b"00000000010001100110101011111010"), -- 1.00795e-38 + -3.61269e-39 = 6.46686e-39
	(b"00000000010101111010011110101111", b"00000000000000000000000000000000"),
	(b"00000000010100000110001111111110", b"00000000101010000000101110101101"), -- 8.04984e-39 + 7.38271e-39 = 1.54326e-38
	(b"10000000001111111010100010101101", b"00000000000000000000000000000000"),
	(b"10000000001111100001100010101101", b"10000000011111011100000101011010"), -- -5.84615e-39 + -5.70265e-39 = -1.15488e-38
	(b"00000000010011100111001010110001", b"00000000000000000000000000000000"),
	(b"10000000011101110110100010001100", b"10000000001010001111010111011011"), -- 7.20431e-39 + -1.09659e-38 = -3.76162e-39
	(b"00000000011000001100100111001000", b"00000000000000000000000000000000"),
	(b"10000000001000100011001110001101", b"00000000001111101001011000111011"), -- 8.88859e-39 + -3.1409e-39 = 5.74769e-39
	(b"00000000000000011110101000000110", b"00000000000000000000000000000000"),
	(b"00000000000111010000101000000101", b"00000000000111101111010000001011"), -- 1.75787e-40 + 2.66682e-39 = 2.84261e-39
	(b"00000000000010111000000110111000", b"00000000000000000000000000000000"),
	(b"00000000000011100000110101010011", b"00000000000110011000111100001011"), -- 1.05672e-39 + 1.29048e-39 = 2.3472e-39
	(b"00000000011001001100110000101101", b"00000000000000000000000000000000"),
	(b"00000000010101001010100011001011", b"00000000101110010111010011111000"), -- 9.25679e-39 + 7.77473e-39 = 1.70315e-38
	(b"00000000010001110100101110010010", b"00000000000000000000000000000000"),
	(b"10000000010000011101000010010110", b"00000000000001010111101011111100"), -- 6.54743e-39 + -6.04413e-39 = 5.03296e-40
	(b"00000000011100111111000011110010", b"00000000000000000000000000000000"),
	(b"10000000000010000101110100110000", b"00000000011010111001001111000010"), -- 1.06475e-38 + -7.68113e-40 = 9.8794e-39
	(b"00000000010110101111101000110000", b"00000000000000000000000000000000"),
	(b"10000000001000011001110010000001", b"00000000001110010101110110101111"), -- 8.35495e-39 + -3.08671e-39 = 5.26823e-39
	(b"00000000001111101000100111000010", b"00000000000000000000000000000000"),
	(b"10000000010111111101100001010110", b"10000000001000010100111010010100"), -- 5.74322e-39 + -8.80198e-39 = -3.05876e-39
	(b"10000000001011110110011010011010", b"00000000000000000000000000000000"),
	(b"10000000010000000100001100000100", b"10000000011011111010100110011110"), -- -4.35307e-39 + -5.90151e-39 = -1.02546e-38
	(b"00000000011101000011011110101100", b"00000000000000000000000000000000"),
	(b"00000000010010000011010011111101", b"00000000101111000110110010101001"), -- 1.06729e-38 + 6.63116e-39 = 1.73041e-38
	(b"00000000001011011110000101111100", b"00000000000000000000000000000000"),
	(b"00000000000100100101011010011100", b"00000000010000000011100000011000"), -- 4.21349e-39 + 1.68411e-39 = 5.89759e-39
	(b"10000000010101011010010010011001", b"00000000000000000000000000000000"),
	(b"10000000010000000100100011001111", b"10000000100101011110110101101000"), -- -7.86506e-39 + -5.90359e-39 = -1.37687e-38
	(b"00000000010110100111000111100001", b"00000000000000000000000000000000"),
	(b"10000000001000000000010011100001", b"00000000001110100110110100000000"), -- 8.30605e-39 + -2.94049e-39 = 5.36556e-39
	(b"00000000000100100011111100110001", b"00000000000000000000000000000000"),
	(b"00000000000000011010100010011011", b"00000000000100111110011111001100"), -- 1.67571e-39 + 1.5232e-40 = 1.82803e-39
	(b"10000000001100101111101001011001", b"00000000000000000000000000000000"),
	(b"00000000000101110010101011010100", b"10000000000110111100111110000101"), -- -4.68158e-39 + 2.12758e-39 = -2.554e-39
	(b"00000000001100101011101110000110", b"00000000000000000000000000000000"),
	(b"10000000011101110011111011010101", b"10000000010001001000001101001111"), -- 4.65905e-39 + -1.0951e-38 = -6.29192e-39
	(b"00000000001100111000000111110010", b"00000000000000000000000000000000"),
	(b"00000000010001100110110010011011", b"00000000011110011110111010001101"), -- 4.73023e-39 + 6.46745e-39 = 1.11977e-38
	(b"10000000000101100000110101000011", b"00000000000000000000000000000000"),
	(b"00000000011001101110111010101110", b"00000000010100001110000101101011"), -- -2.02514e-39 + 9.45284e-39 = 7.4277e-39
	(b"00000000000000011100000110001011", b"00000000000000000000000000000000"),
	(b"00000000000110100001011100100110", b"00000000000110111101100010110001"), -- 1.61266e-40 + 2.39603e-39 = 2.55729e-39
	(b"00000000000111100001101100101111", b"00000000000000000000000000000000"),
	(b"00000000000101100100011001110111", b"00000000001101000110000110100110"), -- 2.76482e-39 + 2.04566e-39 = 4.81048e-39
	(b"10000000000100000001001111010011", b"00000000000000000000000000000000"),
	(b"00000000011100011011101001011100", b"00000000011000011010011010001001"), -- -1.47648e-39 + 1.04443e-38 = 8.96778e-39
	(b"10000000010000011000000011001010", b"00000000000000000000000000000000"),
	(b"00000000001101001111000010010001", b"10000000000011001001000000111001"), -- -6.01551e-39 + 4.86174e-39 = -1.15376e-39
	(b"10000000010110101011111001000100", b"00000000000000000000000000000000"),
	(b"00000000011000101100010001001101", b"00000000000010000000011000001001"), -- -8.33345e-39 + 9.0703e-39 = 7.36849e-40
	(b"00000000010110001101011111000011", b"00000000000000000000000000000000"),
	(b"00000000011110001110010010001101", b"00000000110100011011110001010000"), -- 8.15892e-39 + 1.11022e-38 = 1.92612e-38
	(b"10000000001100010111011110010001", b"00000000000000000000000000000000"),
	(b"00000000000001100010100001011001", b"10000000001010110100111100111000"), -- -4.54283e-39 + 5.65487e-40 = -3.97734e-39
	(b"00000000010101100110111001010010", b"00000000000000000000000000000000"),
	(b"10000000000011011111111110101110", b"00000000010010000110111010100100"), -- 7.93743e-39 + -1.28558e-39 = 6.65185e-39
	(b"00000000000110110101011011111011", b"00000000000000000000000000000000"),
	(b"10000000000110001110001001100111", b"00000000000000100111010010010100"), -- 2.51076e-39 + -2.28527e-39 = 2.25491e-40
	(b"10000000011111100100011011110100", b"00000000000000000000000000000000"),
	(b"10000000001111000101010110111010", b"10000000101110101001110010101110"), -- -1.15967e-38 + -5.54088e-39 = -1.71376e-38
	(b"00000000010101010110011000111001", b"00000000000000000000000000000000"),
	(b"10000000011000010000011110101111", b"10000000000010111010000101110110"), -- 7.84269e-39 + -8.9108e-39 = -1.06811e-39
	(b"00000000001110011100101100011100", b"00000000000000000000000000000000"),
	(b"00000000000001101000000010001000", b"00000000010000000100101110100100"), -- 5.30749e-39 + 5.97121e-40 = 5.90461e-39
	(b"10000000010110111111110001110100", b"00000000000000000000000000000000"),
	(b"00000000001001110011000000100001", b"10000000001101001100110001010011"), -- -8.44759e-39 + 3.59885e-39 = -4.84874e-39
	(b"10000000011000000110001100000001", b"00000000000000000000000000000000"),
	(b"00000000010110110111010010000101", b"10000000000001001110111001111100"), -- -8.85172e-39 + 8.39883e-39 = -4.52894e-40
	(b"00000000001101101011110100010011", b"00000000000000000000000000000000"),
	(b"10000000010001100000001101010111", b"10000000000011110100011001000100"), -- 5.02694e-39 + -6.42968e-39 = -1.40274e-39
	(b"10000000000001101001000001010010", b"00000000000000000000000000000000"),
	(b"00000000000111101011000000000000", b"00000000000110000001111110101110"), -- -6.02785e-40 + 2.8182e-39 = 2.21542e-39
	(b"00000000001010100010001010101100", b"00000000000000000000000000000000"),
	(b"10000000010011011100001100111011", b"10000000001000111010000010001111"), -- 3.86953e-39 + -7.14137e-39 = -3.27184e-39
	(b"00000000011110011100010001100111", b"00000000000000000000000000000000"),
	(b"00000000001011101100011111001001", b"00000000101010001000110000110000"), -- 1.11826e-38 + 4.2961e-39 = 1.54787e-38
	(b"10000000001011000000011001101101", b"00000000000000000000000000000000"),
	(b"00000000000010111001110011111000", b"10000000001000000110100101110101"), -- -4.04307e-39 + 1.0665e-39 = -2.97657e-39
	(b"10000000000110110110100100000101", b"00000000000000000000000000000000"),
	(b"00000000000110011100111100101010", b"10000000000000011001100111011011"), -- -2.51723e-39 + 2.3702e-39 = -1.47028e-40
	(b"10000000001100010000111011111010", b"00000000000000000000000000000000"),
	(b"10000000000101100010101100000010", b"10000000010001110011100111111100"), -- -4.50531e-39 + -2.03581e-39 = -6.54112e-39
	(b"10000000000001011001110011100011", b"00000000000000000000000000000000"),
	(b"10000000011111000010101110111000", b"10000000100000011100100010011011"), -- -5.15458e-40 + -1.14033e-38 = -1.19187e-38
	(b"10000000010101111001000110100110", b"00000000000000000000000000000000"),
	(b"10000000001010101110010110001110", b"10000000100000100111011100110100"), -- -8.04194e-39 + -3.93944e-39 = -1.19814e-38
	(b"10000000001100010110101010110011", b"00000000000000000000000000000000"),
	(b"00000000001001111111111101100110", b"10000000000010010110101101001101"), -- -4.53822e-39 + 3.6732e-39 = -8.65012e-40
	(b"10000000011010010101101100001100", b"00000000000000000000000000000000"),
	(b"10000000011100111111011111010010", b"10000000110111010101001011011110"), -- -9.67539e-39 + -1.065e-38 = -2.03254e-38
	(b"10000000011010111011000110011110", b"00000000000000000000000000000000"),
	(b"00000000000101000100101100101110", b"10000000010101110110011001110000"), -- -9.89012e-39 + 1.86368e-39 = -8.02644e-39
	(b"00000000010101111110100010011000", b"00000000000000000000000000000000"),
	(b"00000000011011100110100100011101", b"00000000110001100101000110110101"), -- 8.07313e-39 + 1.01396e-38 = 1.82127e-38
	(b"00000000001010110101010111010100", b"00000000000000000000000000000000"),
	(b"00000000001001101010001110011001", b"00000000010100011111100101101101"), -- 3.97972e-39 + 3.54844e-39 = 7.52815e-39
	(b"00000000000011100110100101111001", b"00000000000000000000000000000000"),
	(b"10000000001111101001010010110010", b"10000000001100000010101100111001"), -- 1.32353e-39 + -5.74714e-39 = -4.42361e-39
	(b"10000000001101001010001110010011", b"00000000000000000000000000000000"),
	(b"10000000011001000010100101011100", b"10000000100110001100110011101111"), -- -4.83413e-39 + -9.19839e-39 = -1.40325e-38
	(b"10000000010101001000101110001101", b"00000000000000000000000000000000"),
	(b"00000000001010100000011111010111", b"10000000001010101000001110110110"), -- -7.76424e-39 + 3.8599e-39 = -3.90434e-39
	(b"10000000001011010001000100101101", b"00000000000000000000000000000000"),
	(b"00000000000100111100111111101000", b"10000000000110010100000101000101"), -- -4.13876e-39 + 1.81946e-39 = -2.3193e-39
	(b"00000000001011010011010000101100", b"00000000000000000000000000000000"),
	(b"10000000001011011000100001011110", b"10000000000000000101010000110010"), -- 4.15131e-39 + -4.18152e-39 = -3.02036e-41
	(b"00000000011011110101100001100000", b"00000000000000000000000000000000"),
	(b"00000000000111100100010110000101", b"00000000100011011001110111100101"), -- 1.02254e-38 + 2.78e-39 = 1.30054e-38
	(b"10000000010001101101100001001110", b"00000000000000000000000000000000"),
	(b"00000000001110000010110011101000", b"10000000000011101010101101100110"), -- -6.50608e-39 + 5.1589e-39 = -1.34718e-39
	(b"10000000010101101111111011111101", b"00000000000000000000000000000000"),
	(b"00000000011111000010001100111010", b"00000000001001010010010000111101"), -- -7.98933e-39 + 1.14002e-38 = 3.41091e-39
	(b"10000000011001100111101000011111", b"00000000000000000000000000000000"),
	(b"00000000000101010011010111101000", b"10000000010100010100010000110111"), -- -9.41103e-39 + 1.94788e-39 = -7.46315e-39
	(b"00000000011010011011010101001110", b"00000000000000000000000000000000"),
	(b"00000000001000101011000011011011", b"00000000100011000110011000101001"), -- 9.70777e-39 + 3.18585e-39 = 1.28936e-38
	(b"00000000001100011010101101111101", b"00000000000000000000000000000000"),
	(b"10000000001010100010111100110100", b"00000000000001110111110001001001"), -- 4.56146e-39 + -3.87402e-39 = 6.87434e-40
	(b"10000000001011100110100100000010", b"00000000000000000000000000000000"),
	(b"10000000000111111011111000100000", b"10000000010011100010011100100010"), -- -4.2621e-39 + -2.9151e-39 = -7.17721e-39
	(b"10000000000100010110110100010110", b"00000000000000000000000000000000"),
	(b"10000000000010000001101100110001", b"10000000000110011000100001000111"), -- -1.60034e-39 + -7.44438e-40 = -2.34477e-39
	(b"10000000000010101110010000101101", b"00000000000000000000000000000000"),
	(b"10000000000110110101110101100011", b"10000000001001100100000110010000"), -- -1.00021e-39 + -2.51306e-39 = -3.51327e-39
	(b"00000000011000110001001000010000", b"00000000000000000000000000000000"),
	(b"10000000000111111010110001110001", b"00000000010000110110010110011111"), -- 9.09819e-39 + -2.90876e-39 = 6.18943e-39
	(b"00000000000101100000101001010101", b"00000000000000000000000000000000"),
	(b"10000000010101011110000110001111", b"10000000001111111101011100111010"), -- 2.02409e-39 + -7.88693e-39 = -5.86285e-39
	(b"10000000001110000111110011111001", b"00000000000000000000000000000000"),
	(b"00000000001101111001110001100110", b"10000000000000001110000010010011"), -- -5.18762e-39 + 5.10706e-39 = -8.05621e-41
	(b"00000000001011000010111001011011", b"00000000000000000000000000000000"),
	(b"10000000011101111000010000000111", b"10000000010010110101010110101100"), -- 4.05739e-39 + -1.09758e-38 = -6.9184e-39
	(b"00000000011010010001100110000001", b"00000000000000000000000000000000"),
	(b"00000000010001101111010101011101", b"00000000101100000000111011011110"), -- 9.65188e-39 + 6.5165e-39 = 1.61684e-38
	(b"00000000001101100100000110001000", b"00000000000000000000000000000000"),
	(b"00000000001000111110001001010011", b"00000000010110100010001111011011"), -- 4.98262e-39 + 3.29543e-39 = 8.27806e-39
	(b"10000000011011001100000001000100", b"00000000000000000000000000000000"),
	(b"00000000001101000010111001010111", b"10000000001110001001000111101101"), -- -9.98721e-39 + 4.79207e-39 = -5.19514e-39
	(b"00000000010001000111111001001100", b"00000000000000000000000000000000"),
	(b"10000000000000101010111010011011", b"00000000010000011100111110110001"), -- 6.29012e-39 + -2.46308e-40 = 6.04381e-39
	(b"10000000000010001111010011100010", b"00000000000000000000000000000000"),
	(b"10000000011011011110100101000011", b"10000000011101101101111000100101"), -- -8.22531e-40 + -1.00937e-38 = -1.09163e-38
	(b"00000000000100011100110100001110", b"00000000000000000000000000000000"),
	(b"00000000000110101100010000101011", b"00000000001011001001000100111001"), -- 1.63476e-39 + 2.45809e-39 = 4.09286e-39
	(b"00000000011001110100000111101100", b"00000000000000000000000000000000"),
	(b"10000000011100010100101000110001", b"10000000000010100000100001000101"), -- 9.4827e-39 + -1.0404e-38 = -9.21322e-40
	(b"00000000000010100110110100110011", b"00000000000000000000000000000000"),
	(b"10000000000010000101000110101110", b"00000000000000100001101110000101"), -- 9.57528e-40 + -7.63985e-40 = 1.93543e-40
	(b"10000000010000100010100100111110", b"00000000000000000000000000000000"),
	(b"10000000011011110111100011011101", b"10000000101100011010001000011011"), -- -6.07594e-39 + -1.02371e-38 = -1.6313e-38
	(b"10000000010010100001110010011011", b"00000000000000000000000000000000"),
	(b"10000000010000101110011011010110", b"10000000100011010000001101110001"), -- -6.80609e-39 + -6.14395e-39 = -1.295e-38
	(b"10000000000010111110010001011100", b"00000000000000000000000000000000"),
	(b"10000000011111101000011111010001", b"10000000100010100110110000101101"), -- -1.09211e-39 + -1.162e-38 = -1.27121e-38
	(b"00000000001010110110000010101100", b"00000000000000000000000000000000"),
	(b"10000000010100011001111111010011", b"10000000001001100011111100100111"), -- 3.98361e-39 + -7.49601e-39 = -3.5124e-39
	(b"10000000001010011111011110100001", b"00000000000000000000000000000000"),
	(b"10000000001100110011101101101010", b"10000000010111010011001100001011"), -- -3.85409e-39 + -4.70492e-39 = -8.55901e-39
	(b"10000000011100011111010010000100", b"00000000000000000000000000000000"),
	(b"10000000011110011110111000110110", b"10000000111010111110001010111010"), -- -1.04651e-38 + -1.11975e-38 = -2.16627e-38
	(b"10000000000110111101101010001010", b"00000000000000000000000000000000"),
	(b"10000000011001011000101100011101", b"10000000100000010110010110100111"), -- -2.55796e-39 + -9.32529e-39 = -1.18832e-38
	(b"10000000010010111000100001100111", b"00000000000000000000000000000000"),
	(b"10000000001101101101110110000100", b"10000000100000100110010111101011"), -- -6.93659e-39 + -5.03858e-39 = -1.19752e-38
	(b"00000000011100101010001110001101", b"00000000000000000000000000000000"),
	(b"10000000000001010000110000101010", b"00000000011011011001011101100011"), -- 1.05279e-38 + -4.63541e-40 = 1.00644e-38
	(b"00000000001001111101011010010011", b"00000000000000000000000000000000"),
	(b"10000000001110101101000110010110", b"10000000000100101111101100000011"), -- 3.65856e-39 + -5.40164e-39 = -1.74308e-39
	(b"00000000001111101110001100101100", b"00000000000000000000000000000000"),
	(b"10000000011011100101111010111010", b"10000000001011110111101110001110"), -- 5.77529e-39 + -1.01359e-38 = -4.36059e-39
	(b"00000000011110100010101111000101", b"00000000000000000000000000000000"),
	(b"00000000000101100100101101001101", b"00000000100100000111011100010010"), -- 1.12196e-38 + 2.04739e-39 = 1.3267e-38
	(b"00000000001010111110100000010010", b"00000000000000000000000000000000"),
	(b"10000000001000010010111101101001", b"00000000000010101011100010101001"), -- 4.03218e-39 + -3.04758e-39 = 9.84599e-40
	(b"10000000000111111101011011010010", b"00000000000000000000000000000000"),
	(b"00000000011011010110101010010110", b"00000000010011011001001111000100"), -- -2.92396e-39 + 1.00483e-38 = 7.12434e-39
	(b"10000000011111110100111001100100", b"00000000000000000000000000000000"),
	(b"00000000000100011110101100110001", b"10000000011011010110001100110011"), -- -1.16912e-38 + 1.64557e-39 = -1.00457e-38
	(b"00000000011100111101101111010111", b"00000000000000000000000000000000"),
	(b"10000000000110110011010111001011", b"00000000010110001010011000001100"), -- 1.06399e-38 + -2.49886e-39 = 8.14109e-39
	(b"10000000010000100110101101101011", b"00000000000000000000000000000000"),
	(b"10000000001000100111011101101001", b"10000000011001001110001011010100"), -- -6.09968e-39 + -3.16524e-39 = -9.26492e-39
	(b"10000000010111000010010111010001", b"00000000000000000000000000000000"),
	(b"10000000011110100000000110010110", b"10000000110101100010011101100111"), -- -8.46243e-39 + -1.12045e-38 = -1.96669e-38
	(b"10000000000011111110011000100011", b"00000000000000000000000000000000"),
	(b"10000000000110001110010001101101", b"10000000001010001100101010010000"), -- -1.46009e-39 + -2.286e-39 = -3.74609e-39
	(b"10000000001000011011111000010010", b"00000000000000000000000000000000"),
	(b"10000000011110011101100011010000", b"10000000100110111001011011100010"), -- -3.09876e-39 + -1.11899e-38 = -1.42886e-38
	(b"00000000001000000100110010001111", b"00000000000000000000000000000000"),
	(b"10000000011001000100110100101000", b"10000000010001000000000010011001"), -- 2.9662e-39 + -9.21123e-39 = -6.24503e-39
	(b"10000000001001100100110100011100", b"00000000000000000000000000000000"),
	(b"10000000001111110010011010010101", b"10000000011001010111001110110001"), -- -3.51741e-39 + -5.79948e-39 = -9.31689e-39
	(b"10000000011000011100101001000011", b"00000000000000000000000000000000"),
	(b"00000000000010010000101110000111", b"10000000010110001011111010111100"), -- -8.9806e-39 + 8.30655e-40 = -8.14995e-39
	(b"10000000001100101111110000111010", b"00000000000000000000000000000000"),
	(b"10000000000010101010101010001100", b"10000000001111011010011011000110"), -- -4.68226e-39 + -9.79536e-40 = -5.66179e-39
	(b"00000000011010111000101110101011", b"00000000000000000000000000000000"),
	(b"10000000011001011001101111011010", b"00000000000001011110111111010001"), -- 9.8765e-39 + -9.33129e-39 = 5.45207e-40
	(b"10000000001100001010100000000011", b"00000000000000000000000000000000"),
	(b"00000000001000001011110000100100", b"10000000000011111110101111011111"), -- -4.46838e-39 + 3.00623e-39 = -1.46215e-39
	(b"10000000000101100101001101100101", b"00000000000000000000000000000000"),
	(b"10000000001101101110110000011111", b"10000000010011010011111110000100"), -- -2.0503e-39 + -5.04382e-39 = -7.09412e-39
	(b"00000000000111111110001101011001", b"00000000000000000000000000000000"),
	(b"00000000000111101001000000001111", b"00000000001111100111001101101000"), -- 2.92846e-39 + 2.80674e-39 = 5.7352e-39
	(b"10000000001010110100011000000001", b"00000000000000000000000000000000"),
	(b"10000000010100001101011011010101", b"10000000011111000001110011010110"), -- -3.97404e-39 + -7.42391e-39 = -1.13979e-38
	(b"10000000010000110001101100000001", b"00000000000000000000000000000000"),
	(b"10000000000100010001110000001110", b"10000000010101000011011100001111"), -- -6.16267e-39 + -1.57127e-39 = -7.73393e-39
	(b"00000000010001110010001100010001", b"00000000000000000000000000000000"),
	(b"00000000011011001011011110111000", b"00000000101100111101101011001001"), -- 6.5329e-39 + 9.98414e-39 = 1.6517e-38
	(b"00000000010101011000100101110100", b"00000000000000000000000000000000"),
	(b"10000000011010001001111100001001", b"10000000000100110001010110010101"), -- 7.85533e-39 + -9.60794e-39 = -1.75262e-39
	(b"10000000011000100011010000111000", b"00000000000000000000000000000000"),
	(b"00000000011111110101110111111000", b"00000000000111010010100111000000"), -- -9.01861e-39 + 1.16968e-38 = 2.67821e-39
	(b"10000000011111110110110000110000", b"00000000000000000000000000000000"),
	(b"00000000011001110110011000011101", b"10000000000110000000011000010011"), -- -1.17019e-38 + 9.49569e-39 = -2.20623e-39
	(b"10000000010000010111110100010001", b"00000000000000000000000000000000"),
	(b"10000000000010110100100100100000", b"10000000010011001100011000110001"), -- -6.01417e-39 + -1.03642e-39 = -7.0506e-39
	(b"00000000000110011111011001101011", b"00000000000000000000000000000000"),
	(b"00000000001111010000010101001001", b"00000000010101101111101110110100"), -- 2.38429e-39 + 5.60386e-39 = 7.98815e-39
	(b"00000000000100110000000010110110", b"00000000000000000000000000000000"),
	(b"00000000011110000010101111011111", b"00000000100010110010110010010101"), -- 1.74513e-39 + 1.1036e-38 = 1.27811e-38
	(b"00000000010010010110100010011100", b"00000000000000000000000000000000"),
	(b"10000000001001111110001101101000", b"00000000001000011000010100110100"), -- 6.74152e-39 + -3.66316e-39 = 3.07836e-39
	(b"10000000000110111111100100110110", b"00000000000000000000000000000000"),
	(b"00000000000111111101010111000110", b"00000000000000111101110010010000"), -- -2.56896e-39 + 2.92359e-39 = 3.54629e-40
	(b"00000000000111001100111000101010", b"00000000000000000000000000000000"),
	(b"10000000011011101010001110011001", b"10000000010100011101010101101111"), -- 2.64535e-39 + -1.01606e-38 = -7.51524e-39
	(b"00000000011011000101011100101111", b"00000000000000000000000000000000"),
	(b"00000000000100010011011110110000", b"00000000011111011000111011011111"), -- 9.94951e-39 + 1.58118e-39 = 1.15307e-38
	(b"10000000001101101110110100010111", b"00000000000000000000000000000000"),
	(b"00000000010101111110011011111110", b"00000000001000001111100111100111"), -- -5.04417e-39 + 8.07255e-39 = 3.02838e-39
	(b"10000000000100111011011011111101", b"00000000000000000000000000000000"),
	(b"10000000011011011110001111000110", b"10000000100000011001101011000011"), -- -1.81052e-39 + -1.00918e-38 = -1.19023e-38
	(b"10000000001110010011101100101010", b"00000000000000000000000000000000"),
	(b"00000000010111000000101010111001", b"00000000001000101100111110001111"), -- -5.25585e-39 + 8.45271e-39 = 3.19686e-39
	(b"10000000010110101001011011001111", b"00000000000000000000000000000000"),
	(b"10000000000101011100100000111010", b"10000000011100000101111100001001"), -- -8.31929e-39 + -2.00037e-39 = -1.03197e-38
	(b"10000000011100100110100110100000", b"00000000000000000000000000000000"),
	(b"10000000000111001101110011001000", b"10000000100011110100011001101000"), -- -1.05071e-38 + -2.6506e-39 = -1.31577e-38
	(b"00000000011110100011011100000010", b"00000000000000000000000000000000"),
	(b"00000000011001100000000011101101", b"00000000111000000011011111101111"), -- 1.12237e-38 + 9.36755e-39 = 2.05912e-38
	(b"00000000000100001110110011010000", b"00000000000000000000000000000000"),
	(b"10000000000000000111110000101100", b"00000000000100000111000010100100"), -- 1.55432e-39 + -4.45445e-41 = 1.50978e-39
	(b"00000000010100000011100010100011", b"00000000000000000000000000000000"),
	(b"10000000000110111010110110101111", b"00000000001101001000101011110100"), -- 7.36716e-39 + -2.54186e-39 = 4.82529e-39
	(b"00000000001010101111001111000000", b"00000000000000000000000000000000"),
	(b"00000000001001101011101011010100", b"00000000010100011010111010010100"), -- 3.94453e-39 + 3.55677e-39 = 7.5013e-39
	(b"00000000010001101111111000110001", b"00000000000000000000000000000000"),
	(b"00000000001010011101110100111101", b"00000000011100001101101101101110"), -- 6.51967e-39 + 3.84462e-39 = 1.03643e-38
	(b"10000000010011000111111111100000", b"00000000000000000000000000000000"),
	(b"00000000001000111110011101010000", b"10000000001010001001100010010000"), -- -7.02537e-39 + 3.29722e-39 = -3.72815e-39
	(b"00000000011111010010010011110011", b"00000000000000000000000000000000"),
	(b"10000000011010011101111111010010", b"00000000000100110100010100100001"), -- 1.14927e-38 + -9.72302e-39 = 1.76967e-39
	(b"10000000000010001001111100101100", b"00000000000000000000000000000000"),
	(b"10000000011010001000100100000110", b"10000000011100010010100000110010"), -- -7.91784e-40 + -9.60005e-39 = -1.03918e-38
	(b"00000000000001111011111100100100", b"00000000000000000000000000000000"),
	(b"00000000010001010100010011101010", b"00000000010011010000010000001110"), -- 7.11417e-40 + 6.36137e-39 = 7.07279e-39
	(b"00000000000101011100111010100011", b"00000000000000000000000000000000"),
	(b"10000000010111010001011000111001", b"10000000010001110100011110010110"), -- 2.00267e-39 + -8.54867e-39 = -6.546e-39
	(b"10000000010101001111110000010111", b"00000000000000000000000000000000"),
	(b"10000000000010100001101001001011", b"10000000010111110001011001100010"), -- -7.80461e-39 + -9.27787e-40 = -8.7324e-39
	(b"10000000000011100010101111010001", b"00000000000000000000000000000000"),
	(b"10000000011010000110000010100000", b"10000000011101101000110001110001"), -- -1.30142e-39 + -9.58555e-39 = -1.0887e-38
	(b"10000000001101010001000001101110", b"00000000000000000000000000000000"),
	(b"10000000000100001111100000001010", b"10000000010001100000100001111000"), -- -4.87318e-39 + -1.55835e-39 = -6.43152e-39
	(b"00000000010101011001001000011101", b"00000000000000000000000000000000"),
	(b"10000000010011000001000011111110", b"00000000000010011000000100011111"), -- 7.85843e-39 + -6.98559e-39 = 8.72839e-40
	(b"10000000000110000010110100011111", b"00000000000000000000000000000000"),
	(b"10000000001000111010101001001000", b"10000000001110111101011101100111"), -- -2.22024e-39 + -3.27533e-39 = -5.49557e-39
	(b"00000000000100100001110000001011", b"00000000000000000000000000000000"),
	(b"00000000011101110000001011000101", b"00000000100010010001111011010000"), -- 1.6631e-39 + 1.09294e-38 = 1.25925e-38
	(b"00000000011111010101001010111111", b"00000000000000000000000000000000"),
	(b"10000000010000110010111111000110", b"00000000001110100010001011111001"), -- 1.15091e-38 + -6.17012e-39 = 5.339e-39
	(b"00000000011010110001001111110101", b"00000000000000000000000000000000"),
	(b"00000000011101001010011000000111", b"00000000110111111011100111111100"), -- 9.83356e-39 + 1.07125e-38 = 2.0546e-38
	(b"10000000001011101010111101101100", b"00000000000000000000000000000000"),
	(b"10000000011100000100111001010010", b"10000000100111101111110110111110"), -- -4.28736e-39 + -1.03137e-38 = -1.4601e-38
	(b"00000000000001001100011011101010", b"00000000000000000000000000000000"),
	(b"00000000000001000011101011000101", b"00000000000010010000000110101111"), -- 4.38699e-40 + 3.88425e-40 = 8.27123e-40
	(b"10000000011001000001001111110101", b"00000000000000000000000000000000"),
	(b"10000000001111010101011010010110", b"10000000101000010110101010001011"), -- -9.19071e-39 + -5.63303e-39 = -1.48237e-38
	(b"00000000001011000101101111110111", b"00000000000000000000000000000000"),
	(b"10000000011010100100111100011110", b"10000000001111011111001100100111"), -- 4.07375e-39 + -9.76294e-39 = -5.68919e-39
	(b"00000000010101111111010010000111", b"00000000000000000000000000000000"),
	(b"00000000001001101001101010111100", b"00000000011111101000111101000011"), -- 8.07741e-39 + 3.54526e-39 = 1.16227e-38
	(b"00000000011101101001111010001101", b"00000000000000000000000000000000"),
	(b"10000000001111111000001010010001", b"00000000001101110001101111111100"), -- 1.08935e-38 + -5.83247e-39 = 5.06099e-39
	(b"10000000011001100011010010010010", b"00000000000000000000000000000000"),
	(b"00000000001100000001110010110110", b"10000000001101100001011111011100"), -- -9.38608e-39 + 4.4184e-39 = -4.96768e-39
	(b"10000000000111011011011110110101", b"00000000000000000000000000000000"),
	(b"10000000001110000100011011010110", b"10000000010101011111111010001011"), -- -2.72913e-39 + -5.1682e-39 = -7.89733e-39
	(b"00000000000001110010010010100000", b"00000000000000000000000000000000"),
	(b"10000000010001110110000101000011", b"10000000010000000011110010100011"), -- 6.55987e-40 + -6.55521e-39 = -5.89922e-39
	(b"10000000001001010111111011010101", b"00000000000000000000000000000000"),
	(b"00000000001101111001110111011110", b"00000000000100100001111100001001"), -- -3.44341e-39 + 5.10758e-39 = 1.66417e-39
	(b"00000000011000010101101111010111", b"00000000000000000000000000000000"),
	(b"10000000000011111001100000110101", b"00000000010100011100001110100010"), -- 8.94099e-39 + -1.43213e-39 = 7.50886e-39
	(b"10000000001110010011100111111000", b"00000000000000000000000000000000"),
	(b"00000000011110000111100111110111", b"00000000001111110011111111111111"), -- -5.25542e-39 + 1.1064e-38 = 5.80859e-39
	(b"00000000001011000001100110010010", b"00000000000000000000000000000000"),
	(b"10000000010100000100110111010000", b"10000000001001000011010000111110"), -- 4.04993e-39 + -7.37475e-39 = -3.32482e-39
	(b"10000000000010101011101010111110", b"00000000000000000000000000000000"),
	(b"10000000001100100100000011001110", b"10000000001111001111101110001100"), -- -9.85345e-40 + -4.61502e-39 = -5.60037e-39
	(b"10000000010111110111101000011111", b"00000000000000000000000000000000"),
	(b"10000000001001100111000110010010", b"10000000100001011110101110110001"), -- -8.76818e-39 + -3.53049e-39 = -1.22987e-38
	(b"00000000000101011111100011101111", b"00000000000000000000000000000000"),
	(b"00000000010010100101001010000100", b"00000000011000000100101101110011"), -- 2.01785e-39 + 6.82543e-39 = 8.84327e-39
	(b"00000000000101101100100001111111", b"00000000000000000000000000000000"),
	(b"00000000001001010010111110101110", b"00000000001110111111100000101101"), -- 2.09231e-39 + 3.41502e-39 = 5.50732e-39
	(b"00000000010101010100111010110001", b"00000000000000000000000000000000"),
	(b"10000000011000011011101000110111", b"10000000000011000110101110000110"), -- 7.83425e-39 + -8.97484e-39 = -1.1406e-39
	(b"10000000010111101101010100111111", b"00000000000000000000000000000000"),
	(b"00000000000010000100101110000000", b"10000000010101101000100110111111"), -- -8.70903e-39 + 7.61768e-40 = -7.94727e-39
	(b"10000000001100001100111110001011", b"00000000000000000000000000000000"),
	(b"00000000011010011010111101011111", b"00000000001110001101111111010100"), -- -4.48256e-39 + 9.70564e-39 = 5.22308e-39
	(b"00000000001111011101100110110000", b"00000000000000000000000000000000"),
	(b"00000000011100110110010101101101", b"00000000101100010011111100011101"), -- 5.68006e-39 + 1.05975e-38 = 1.62775e-38
	(b"10000000001000100101110000111111", b"00000000000000000000000000000000"),
	(b"00000000000010000111101110001011", b"10000000000110011110000010110100"), -- -3.1555e-39 + 7.79003e-40 = -2.3765e-39
	(b"10000000001011101101110101100001", b"00000000000000000000000000000000"),
	(b"00000000001101100111110111100011", b"00000000000001111010000010000010"), -- -4.30385e-39 + 5.00428e-39 = 7.00428e-40
	(b"00000000000011111110100100000000", b"00000000000000000000000000000000"),
	(b"00000000011100101101110101011101", b"00000000100000101100011001011101"), -- 1.46112e-39 + 1.05487e-38 = 1.20098e-38
	(b"10000000010101011101101101000111", b"00000000000000000000000000000000"),
	(b"00000000001001000001100011101001", b"10000000001100011100001001011110"), -- -7.88468e-39 + 3.31501e-39 = -4.56967e-39
	(b"10000000010101000001010000101001", b"00000000000000000000000000000000"),
	(b"00000000000011101000110000000111", b"10000000010001011000100000100010"), -- -7.72141e-39 + 1.33593e-39 = -6.38548e-39
	(b"00000000010111010111101100101101", b"00000000000000000000000000000000"),
	(b"10000000011011100010110101100101", b"10000000000100001011001000111000"), -- 8.58489e-39 + -1.01182e-38 = -1.5333e-39
	(b"10000000010100110010000101110010", b"00000000000000000000000000000000"),
	(b"10000000010011100001101101000001", b"10000000101000010011110010110011"), -- -7.63434e-39 + -7.17295e-39 = -1.48073e-38
	(b"10000000001110101010111101000000", b"00000000000000000000000000000000"),
	(b"00000000001110001110000101001010", b"10000000000000011100110111110110"), -- -5.38933e-39 + 5.22361e-39 = -1.6572e-40
	(b"00000000011101101110101111111110", b"00000000000000000000000000000000"),
	(b"10000000011111001101110100010101", b"10000000000001011111000100010111"), -- 1.09212e-38 + -1.14669e-38 = -5.45664e-40
	(b"00000000000100010001000111100101", b"00000000000000000000000000000000"),
	(b"00000000011001011101010110111000", b"00000000011101101110011110011101"), -- 1.56762e-39 + 9.35205e-39 = 1.09197e-38
	(b"10000000000000001001111011001110", b"00000000000000000000000000000000"),
	(b"00000000000111111000011111100110", b"00000000000111101110100100011000"), -- -5.69684e-41 + 2.89565e-39 = 2.83868e-39
	(b"00000000011101101101100001010100", b"00000000000000000000000000000000"),
	(b"00000000010100010001000011000010", b"00000000110001111110100100010110"), -- 1.09142e-38 + 7.44469e-39 = 1.83589e-38
	(b"00000000010010010010011101011100", b"00000000000000000000000000000000"),
	(b"10000000000001100111100101000010", b"00000000010000101010111000011010"), -- 6.71811e-39 + -5.94512e-40 = 6.1236e-39
	(b"00000000000000101100010000111110", b"00000000000000000000000000000000"),
	(b"10000000000101010110110101111011", b"10000000000100101010100100111101"), -- 2.54069e-40 + -1.96782e-39 = -1.71375e-39
	(b"00000000010010001110010100000110", b"00000000000000000000000000000000"),
	(b"00000000010011101101010110100100", b"00000000100101111011101010101010"), -- 6.69431e-39 + 7.23981e-39 = 1.39341e-38
	(b"10000000010101001101110100001100", b"00000000000000000000000000000000"),
	(b"10000000010101000001011110001000", b"10000000101010001111010010010100"), -- -7.79348e-39 + -7.72262e-39 = -1.55161e-38
	(b"10000000010100011110101100001011", b"00000000000000000000000000000000"),
	(b"10000000010111101010000111011011", b"10000000101100001000110011100110"), -- -7.52299e-39 + -8.6906e-39 = -1.62136e-38
	(b"00000000010001100111100011111101", b"00000000000000000000000000000000"),
	(b"00000000000010000011000100010011", b"00000000010011101010101000010000"), -- 6.47189e-39 + 7.52288e-40 = 7.22418e-39
	(b"10000000001101011000011111100100", b"00000000000000000000000000000000"),
	(b"00000000001100101010100111100100", b"10000000000000101101111000000000"), -- -4.91603e-39 + 4.65272e-39 = -2.6331e-40
	(b"10000000010001001001110101000001", b"00000000000000000000000000000000"),
	(b"10000000011110101111001011101110", b"10000000101111111001000000101111"), -- -6.30123e-39 + -1.12911e-38 = -1.75923e-38
	(b"10000000001101011100100100110100", b"00000000000000000000000000000000"),
	(b"10000000010101111010100100100110", b"10000000100011010111001001011010"), -- -4.93946e-39 + -8.05037e-39 = -1.29898e-38
	(b"10000000000001101000110011100010", b"00000000000000000000000000000000"),
	(b"00000000000101100011110011111010", b"00000000000011111011000000011000"), -- -6.01552e-40 + 2.04226e-39 = 1.4407e-39
	(b"10000000010010000111110111110011", b"00000000000000000000000000000000"),
	(b"10000000010010010110110010010101", b"10000000100100011110101010001000"), -- -6.65734e-39 + -6.74294e-39 = -1.34003e-38
	(b"10000000011010011101010001010011", b"00000000000000000000000000000000"),
	(b"00000000000111100111011011111100", b"10000000010010110101110101010111"), -- -9.71889e-39 + 2.79775e-39 = -6.92115e-39
	(b"00000000000100100101000011001000", b"00000000000000000000000000000000"),
	(b"10000000010001100100100101001010", b"10000000001100111111100010000010"), -- 1.68202e-39 + -6.45478e-39 = -4.77276e-39
	(b"00000000010100001011100001000000", b"00000000000000000000000000000000"),
	(b"00000000011001100101100000110001", b"00000000101101110001000001110001"), -- 7.41294e-39 + 9.39886e-39 = 1.68118e-38
	(b"00000000010110010111001100001001", b"00000000000000000000000000000000"),
	(b"00000000000000101000100111001010", b"00000000010110111111110011010011"), -- 8.21463e-39 + 2.331e-40 = 8.44773e-39
	(b"00000000011011010111111001011111", b"00000000000000000000000000000000"),
	(b"00000000010001011111100101110011", b"00000000101100110111011111010010"), -- 1.00554e-38 + 6.42613e-39 = 1.64815e-38
	(b"10000000000000011011111110100100", b"00000000000000000000000000000000"),
	(b"00000000010001010111010011101000", b"00000000010000111011010101000100"), -- -1.60583e-40 + 6.37859e-39 = 6.218e-39
	(b"10000000000100101101110001011011", b"00000000000000000000000000000000"),
	(b"00000000011010011101000100110011", b"00000000010101101111010011011000"), -- -1.73209e-39 + 9.71777e-39 = 7.98569e-39
	(b"00000000001101010101001101110010", b"00000000000000000000000000000000"),
	(b"10000000001100110000100110010001", b"00000000000000100100100111100001"), -- 4.89722e-39 + -4.68704e-39 = 2.10174e-40
	(b"00000000010100111111101110010111", b"00000000000000000000000000000000"),
	(b"10000000011000110110001000001001", b"10000000000011110110011001110010"), -- 7.7126e-39 + -9.12688e-39 = -1.41428e-39
	(b"00000000000101001110001000101100", b"00000000000000000000000000000000"),
	(b"00000000000011110100000000101101", b"00000000001001000010001001011001"), -- 1.91785e-39 + 1.40055e-39 = 3.3184e-39
	(b"10000000010110011110011111110101", b"00000000000000000000000000000000"),
	(b"10000000001101101001110010010100", b"10000000100100001000010010001001"), -- -8.25657e-39 + -5.01529e-39 = -1.32719e-38
	(b"00000000011110101001111111001101", b"00000000000000000000000000000000"),
	(b"00000000010000101010011010101010", b"00000000101111010100011001110111"), -- 1.12613e-38 + 6.12093e-39 = 1.73822e-38
	(b"00000000001111000101101101111100", b"00000000000000000000000000000000"),
	(b"00000000010000001110111110101111", b"00000000011111010100101100101011"), -- 5.54295e-39 + 5.96345e-39 = 1.15064e-38
	(b"10000000010101101010000100101100", b"00000000000000000000000000000000"),
	(b"00000000011110011111010001011111", b"00000000001000110101001100110011"), -- -7.95567e-39 + 1.11998e-38 = 3.24409e-39
	(b"10000000000000011001010111001010", b"00000000000000000000000000000000"),
	(b"10000000000011111010110010000001", b"10000000000100010100001001001011"), -- -1.4557e-40 + -1.43942e-39 = -1.58498e-39
	(b"10000000000001000011010111000011", b"00000000000000000000000000000000"),
	(b"00000000010100111011110011010101", b"00000000010011111000011100010010"), -- -3.86628e-40 + 7.69009e-39 = 7.30346e-39
	(b"10000000000010100111011000111001", b"00000000000000000000000000000000"),
	(b"00000000010101001001110010001110", b"00000000010010100010011001010101"), -- -9.60765e-40 + 7.77034e-39 = 6.80958e-39
	(b"00000000001100000001111100011111", b"00000000000000000000000000000000"),
	(b"10000000000010100110000100010010", b"00000000001001011011111000001101"), -- 4.41927e-39 + -9.53177e-40 = 3.46609e-39
	(b"00000000001110111001001000010100", b"00000000000000000000000000000000"),
	(b"10000000011000111110011111011100", b"10000000001010000101010111001000"), -- 5.4707e-39 + -9.17489e-39 = -3.70419e-39
	(b"00000000010011101100110111110100", b"00000000000000000000000000000000"),
	(b"00000000001000111001000101100001", b"00000000011100100101111101010101"), -- 7.23705e-39 + 3.26639e-39 = 1.05034e-38
	(b"10000000000101111111110011111110", b"00000000000000000000000000000000"),
	(b"00000000010111110111100000100100", b"00000000010001110111101100100110"), -- -2.20297e-39 + 8.76747e-39 = 6.5645e-39
	(b"00000000010000000110100110111110", b"00000000000000000000000000000000"),
	(b"10000000001111001110100110000100", b"00000000000000111000000000111010"), -- 5.9154e-39 + -5.5939e-39 = 3.21506e-40
	(b"00000000000111111011011001100101", b"00000000000000000000000000000000"),
	(b"00000000000011100100011100110110", b"00000000001011011111110110011011"), -- 2.91233e-39 + 1.31124e-39 = 4.22357e-39
	(b"00000000001011101101010110011110", b"00000000000000000000000000000000"),
	(b"10000000010101111111100100001011", b"10000000001010010010001101101101"), -- 4.30106e-39 + -8.07903e-39 = -3.77796e-39
	(b"00000000001111001110001010110010", b"00000000000000000000000000000000"),
	(b"00000000001001100001000110101110", b"00000000011000101111010001100000"), -- 5.59145e-39 + 3.49609e-39 = 9.08754e-39
	(b"00000000001100100101101011010111", b"00000000000000000000000000000000"),
	(b"00000000010111011010010101111011", b"00000000100100000000000001010010"), -- 4.62436e-39 + 8.60006e-39 = 1.32244e-38
	(b"10000000010100011001101000011001", b"00000000000000000000000000000000"),
	(b"10000000010110100110101001100010", b"10000000101011000000010001111011"), -- -7.49396e-39 + -8.30336e-39 = -1.57973e-38
	(b"00000000010100001011010010100100", b"00000000000000000000000000000000"),
	(b"10000000010111101001100110101011", b"10000000000011011110010100000111"), -- 7.41164e-39 + -8.68766e-39 = -1.27602e-39
	(b"10000000010101001011000011100100", b"00000000000000000000000000000000"),
	(b"00000000010111110001001111111010", b"00000000000010100110001100010110"), -- -7.77764e-39 + 8.73154e-39 = 9.539e-40
	(b"10000000001000101101000111011100", b"00000000000000000000000000000000"),
	(b"00000000011101100111000110010000", b"00000000010100111001111110110100"), -- -3.19769e-39 + 1.08773e-38 = 7.67964e-39
	(b"00000000011011101110100111101001", b"00000000000000000000000000000000"),
	(b"00000000000100100000110011000001", b"00000000100000001111011010101010"), -- 1.01858e-38 + 1.65761e-39 = 1.18434e-38
	(b"00000000011101010111001001100100", b"00000000000000000000000000000000"),
	(b"00000000010111110010111100010000", b"00000000110101001010000101110100"), -- 1.07858e-38 + 8.74125e-39 = 1.9527e-38
	(b"10000000010111011100110100101111", b"00000000000000000000000000000000"),
	(b"10000000010011111010000110000101", b"10000000101011010110111010110100"), -- -8.61431e-39 + -7.31295e-39 = -1.59273e-38
	(b"00000000011101010100010011100110", b"00000000000000000000000000000000"),
	(b"10000000001100110010101010110011", b"00000000010000100001101000110011"), -- 1.07695e-38 + -4.69893e-39 = 6.07054e-39
	(b"10000000010100011001000010100000", b"00000000000000000000000000000000"),
	(b"00000000011011011100100100011100", b"00000000000111000011100001111100"), -- -7.49056e-39 + 1.00822e-38 = 2.59166e-39
	(b"00000000011111000111001001111010", b"00000000000000000000000000000000"),
	(b"00000000000011011101100101101011", b"00000000100010100100101111100101"), -- 1.14287e-38 + 1.27186e-39 = 1.27005e-38
	(b"00000000011000101000011001011001", b"00000000000000000000000000000000"),
	(b"10000000000011010110001100111101", b"00000000010101010010001100011100"), -- 9.04807e-39 + -1.22946e-39 = 7.81861e-39
	(b"00000000011110110101110011100001", b"00000000000000000000000000000000"),
	(b"10000000010000000010111000011010", b"00000000001110110010111011000111"), -- 1.13291e-38 + -5.89401e-39 = 5.43507e-39
	(b"10000000000001011010000000000000", b"00000000000000000000000000000000"),
	(b"00000000011011100000011101011101", b"00000000011010000110011101011101"), -- -5.16575e-40 + 1.01045e-38 = 9.58797e-39
	(b"00000000000100001111100001010010", b"00000000000000000000000000000000"),
	(b"00000000010100100111111111001001", b"00000000011000110111100000011011"), -- 1.55845e-39 + 7.57635e-39 = 9.1348e-39
	(b"10000000000100010010101110010100", b"00000000000000000000000000000000"),
	(b"00000000010100110100011101000110", b"00000000010000100001101110110010"), -- -1.57684e-39 + 7.64791e-39 = 6.07108e-39
	(b"00000000000011010101101100011110", b"00000000000000000000000000000000"),
	(b"10000000010100001100100010101011", b"10000000010000110110110110001101"), -- 1.22655e-39 + -7.41883e-39 = -6.19228e-39
	(b"00000000011110011010011110101100", b"00000000000000000000000000000000"),
	(b"10000000011001110110010000001010", b"00000000000100100100001110100010"), -- 1.11722e-38 + -9.49494e-39 = 1.6773e-39
	(b"10000000000100111000011000011010", b"00000000000000000000000000000000"),
	(b"00000000011001110010100000001011", b"00000000010100111010000111110001"), -- -1.79298e-39 + 9.47342e-39 = 7.68044e-39
	(b"10000000000010100110110000001010", b"00000000000000000000000000000000"),
	(b"10000000011010001101010111110011", b"10000000011100110100000111111101"), -- -9.57112e-40 + -9.62764e-39 = -1.05848e-38
	(b"10000000011101101000011000001011", b"00000000000000000000000000000000"),
	(b"00000000001100111000100101001000", b"10000000010000101111110011000011"), -- -1.08847e-38 + 4.73286e-39 = -6.15182e-39
	(b"00000000010111111110100010000010", b"00000000000000000000000000000000"),
	(b"10000000010010001111001101010010", b"00000000000101101111010100110000"), -- 8.80778e-39 + -6.69944e-39 = 2.10834e-39
	(b"10000000010011010101011010001111", b"00000000000000000000000000000000"),
	(b"00000000010010000000001111110100", b"10000000000001010101001010011011"), -- -7.10238e-39 + 6.61357e-39 = -4.88811e-40
	(b"10000000011100000100100111101111", b"00000000000000000000000000000000"),
	(b"10000000011110110011000000011010", b"10000000111010110111101000001001"), -- -1.03121e-38 + -1.1313e-38 = -2.16251e-38
	(b"00000000000001001010000110010011", b"00000000000000000000000000000000"),
	(b"00000000000111001101001100001110", b"00000000001000010111010010100001"), -- 4.25304e-40 + 2.64711e-39 = 3.07241e-39
	(b"00000000001101011001001110010011", b"00000000000000000000000000000000"),
	(b"00000000000000101101110000110010", b"00000000001110000110111111000101"), -- 4.92022e-39 + 2.62662e-40 = 5.18288e-39
	(b"10000000000001111111110100100101", b"00000000000000000000000000000000"),
	(b"10000000000111011011100011011011", b"10000000001001011011011000000000"), -- -7.3366e-40 + -2.72954e-39 = -3.4632e-39
	(b"10000000000100011001111010000010", b"00000000000000000000000000000000"),
	(b"00000000011101100100110001010001", b"00000000011001001010110111001111"), -- -1.61807e-39 + 1.0864e-38 = 9.2459e-39
	(b"00000000010010001010110101011111", b"00000000000000000000000000000000"),
	(b"10000000001000111011011001011011", b"00000000001001001111011100000100"), -- 6.67435e-39 + -3.27966e-39 = 3.39469e-39
	(b"00000000000010101001011110000000", b"00000000000000000000000000000000"),
	(b"10000000000000101100101111110110", b"00000000000001111100101110001010"), -- 9.72703e-40 + -2.56838e-40 = 7.15865e-40
	(b"10000000011100101001100001111100", b"00000000000000000000000000000000"),
	(b"10000000000101001111111100111000", b"10000000100001111001011110110100"), -- -1.05239e-38 + -1.92827e-39 = -1.24522e-38
	(b"10000000011000001100111101111010", b"00000000000000000000000000000000"),
	(b"10000000010011101101000001110110", b"10000000101011111001111111110000"), -- -8.89064e-39 + -7.23795e-39 = -1.61286e-38
	(b"00000000000010100101000100100001", b"00000000000000000000000000000000"),
	(b"00000000001101000001110110001010", b"00000000001111100110111010101011"), -- 9.47459e-40 + 4.78604e-39 = 5.7335e-39
	(b"00000000010011111010010111100100", b"00000000000000000000000000000000"),
	(b"00000000010100011011000111110000", b"00000000101000010101011111010100"), -- 7.31451e-39 + 7.50251e-39 = 1.4817e-38
	(b"00000000010011010111110101000010", b"00000000000000000000000000000000"),
	(b"10000000010111111101100000110110", b"10000000000100100101101011110100"), -- 7.11627e-39 + -8.80193e-39 = -1.68567e-39
	(b"00000000011001101111101100000011", b"00000000000000000000000000000000"),
	(b"00000000011010111001011100101011", b"00000000110100101001001000101110"), -- 9.45727e-39 + 9.88063e-39 = 1.93379e-38
	(b"10000000001001010111001100011011", b"00000000000000000000000000000000"),
	(b"00000000010110110110100110100000", b"00000000001101011111011010000101"), -- -3.43921e-39 + 8.39492e-39 = 4.95572e-39
	(b"10000000001101010110100100111011", b"00000000000000000000000000000000"),
	(b"00000000001101010011011111111000", b"10000000000000000011000101000011"), -- -4.90503e-39 + 4.88736e-39 = -1.76718e-41
	(b"10000000010000100111011000011111", b"00000000000000000000000000000000"),
	(b"10000000010110011100000101100101", b"10000000100111000011011110000100"), -- -6.10352e-39 + -8.24274e-39 = -1.43463e-38
	(b"00000000001110101101110110100111", b"00000000000000000000000000000000"),
	(b"00000000000010101010011011001111", b"00000000010001011000010001110110"), -- 5.40597e-39 + 9.78195e-40 = 6.38417e-39
	(b"10000000010110000110000111011011", b"00000000000000000000000000000000"),
	(b"10000000010101111011101111000101", b"10000000101100000001110110100000"), -- -8.11663e-39 + -8.05705e-39 = -1.61737e-38
	(b"00000000011011111111100101111100", b"00000000000000000000000000000000"),
	(b"00000000011001010101000101111111", b"00000000110101010100101011111011"), -- 1.02832e-38 + 9.30462e-39 = 1.95879e-38
	(b"00000000001011011110011010110010", b"00000000000000000000000000000000"),
	(b"10000000010100100100011101011001", b"10000000001001000110000010100111"), -- 4.21536e-39 + -7.55611e-39 = -3.34075e-39
	(b"00000000011011000100011010000000", b"00000000000000000000000000000000"),
	(b"10000000010010011100001010100000", b"00000000001000101000001111100000"), -- 9.94352e-39 + -6.77381e-39 = 3.16971e-39
	(b"00000000000110000101111111101000", b"00000000000000000000000000000000"),
	(b"00000000001010011100011011011110", b"00000000010000100010011011000110"), -- 2.23846e-39 + 3.8366e-39 = 6.07505e-39
	(b"10000000010011110001110011010100", b"00000000000000000000000000000000"),
	(b"10000000011001100000000100101110", b"10000000101101010001111000000010"), -- -7.26535e-39 + -9.36764e-39 = -1.6633e-38
	(b"00000000011000101101010000111100", b"00000000000000000000000000000000"),
	(b"00000000010000110011011001011100", b"00000000101001100000101010011000"), -- 9.07601e-39 + 6.17248e-39 = 1.52485e-38
	(b"00000000011101110001111010100100", b"00000000000000000000000000000000"),
	(b"00000000011011011110001001010000", b"00000000111001010000000011110100"), -- 1.09394e-38 + 1.00913e-38 = 2.10307e-38
	(b"10000000011100101011101001001000", b"00000000000000000000000000000000"),
	(b"10000000011110111000101101101101", b"10000000111011100100010110110101"), -- -1.05361e-38 + -1.13458e-38 = -2.18819e-38
	(b"10000000000101111011001100000101", b"00000000000000000000000000000000"),
	(b"00000000000010000000011001111101", b"10000000000011111010110010001000"), -- -2.17644e-39 + 7.37012e-40 = -1.43942e-39
	(b"10000000010010000101011000010011", b"00000000000000000000000000000000"),
	(b"00000000001100111100011011100010", b"10000000000101001000111100110001"), -- -6.64303e-39 + 4.75496e-39 = -1.88808e-39
	
	(b"10000000001001010110001010100101", b"00000000000000000000000000000000"),
	(b"10000000010011000000000110101110", b"10000000011100010110010001010011"), -- -3.4333e-39 + -6.9801e-39 = -1.04134e-38
	(b"00000000011001100110110110010111", b"00000000000000000000000000000000"),
	(b"10000000011111101100001101100011", b"10000000000110000101010111001100"), -- 9.40653e-39 + -1.16414e-38 = -2.23483e-39
	(b"00000000000100001011001011111101", b"00000000000000000000000000000000"),
	(b"10000000001001111011110000110101", b"10000000000101110000100100111000"), -- 1.53358e-39 + -3.6491e-39 = -2.11552e-39
	(b"10000000010101001101111000110010", b"00000000000000000000000000000000"),
	(b"10000000011011101100000111101111", b"10000000110000111010000000100001"), -- -7.79389e-39 + -1.01715e-38 = -1.79654e-38
	(b"10000000001101100000001011010101", b"00000000000000000000000000000000"),
	(b"00000000010111110010001010100001", b"00000000001010010001111111001100"), -- -4.96013e-39 + 8.73679e-39 = 3.77666e-39
	(b"00000000010010000001011101100100", b"00000000000000000000000000000000"),
	(b"10000000000101001101001110001011", b"00000000001100110100001111011001"), -- 6.62055e-39 + -1.9126e-39 = 4.70795e-39
	(b"10000000000111000110010111111100", b"00000000000000000000000000000000"),
	(b"00000000010111001010100001111000", b"00000000010000000100001001111100"), -- -2.60798e-39 + 8.5093e-39 = 5.90132e-39
	(b"00000000011100110000101101101110", b"00000000000000000000000000000000"),
	(b"00000000011110011100100111001101", b"00000000111011001101010100111011"), -- 1.05652e-38 + 1.11845e-38 = 2.17497e-38
	(b"10000000001100000101010100001001", b"00000000000000000000000000000000"),
	(b"10000000000000011010001010100000", b"10000000001100011111011110101001"), -- -4.43861e-39 + -1.50174e-40 = -4.58878e-39
	(b"00000000011100000010100010011110", b"00000000000000000000000000000000"),
	(b"10000000010000101110011001110001", b"00000000001011010100001000101101"), -- 1.03001e-38 + -6.14381e-39 = 4.15634e-39
	(b"00000000010100101110000001100010", b"00000000000000000000000000000000"),
	(b"00000000010101001000101111100001", b"00000000101001110110110001000011"), -- 7.611e-39 + 7.76436e-39 = 1.53754e-38
	(b"10000000000001000100000011000010", b"00000000000000000000000000000000"),
	(b"10000000001110010001010100011000", b"10000000001111010101010111011010"), -- -3.90573e-40 + -5.24219e-39 = -5.63276e-39
	(b"00000000010110001010000100000111", b"00000000000000000000000000000000"),
	(b"10000000001111100001100101101001", b"00000000000110101000011110011110"), -- 8.13929e-39 + -5.70292e-39 = 2.43637e-39
	(b"10000000000110000101001111000001", b"00000000000000000000000000000000"),
	(b"10000000001010001101001110110001", b"10000000010000010010011101110010"), -- -2.2341e-39 + -3.74936e-39 = -5.98346e-39
	(b"00000000010010010110110001011000", b"00000000000000000000000000000000"),
	(b"10000000000001010001010110010100", b"00000000010001000101011011000100"), -- 6.74286e-39 + -4.66918e-40 = 6.27594e-39
	(b"10000000010010101100000111010000", b"00000000000000000000000000000000"),
	(b"00000000000011111001010111100001", b"10000000001110110010101111101111"), -- -6.86535e-39 + 1.4313e-39 = -5.43405e-39
	(b"00000000010101000100110101111001", b"00000000000000000000000000000000"),
	(b"10000000001100010100011000110001", b"00000000001000110000011101001000"), -- 7.74197e-39 + -4.52512e-39 = 3.21685e-39
	(b"10000000001100010010010110110101", b"00000000000000000000000000000000"),
	(b"10000000011011111000000111010100", b"10000000101000001010011110001001"), -- -4.51347e-39 + -1.02403e-38 = -1.47538e-38
	(b"00000000001000011100001011101000", b"00000000000000000000000000000000"),
	(b"00000000000001100111001110010001", b"00000000001010000011011001111001"), -- 3.10049e-39 + 5.9247e-40 = 3.69296e-39
	(b"10000000000001101000010011100111", b"00000000000000000000000000000000"),
	(b"10000000011111011100100100001001", b"10000000100001000100110111110000"), -- -5.98689e-40 + -1.15516e-38 = -1.21502e-38
	(b"00000000000011010110010111100101", b"00000000000000000000000000000000"),
	(b"10000000011111001010100111001011", b"10000000011011110100001111100110"), -- 1.23041e-39 + -1.14485e-38 = -1.02181e-38
	(b"10000000001001000010001001011101", b"00000000000000000000000000000000"),
	(b"10000000010111111110010001001101", b"10000000100001000000011010101010"), -- -3.31841e-39 + -8.80627e-39 = -1.21247e-38
	(b"00000000010110010100010100101100", b"00000000000000000000000000000000"),
	(b"10000000011101010011101010101011", b"10000000000110111111010101111111"), -- 8.19817e-39 + -1.07658e-38 = -2.56763e-39
	(b"10000000011001110001111101110110", b"00000000000000000000000000000000"),
	(b"10000000001111101000101100001001", b"10000000101001011010101001111111"), -- -9.47034e-39 + -5.74368e-39 = -1.5214e-38
	(b"00000000010100010011110110010110", b"00000000000000000000000000000000"),
	(b"00000000011001111011100111110011", b"00000000101110001111011110001001"), -- 7.46077e-39 + 9.52576e-39 = 1.69865e-38
	(b"10000000011111000010011101010000", b"00000000000000000000000000000000"),
	(b"10000000001100101001100011101111", b"10000000101011101100000000111111"), -- -1.14017e-38 + -4.64664e-39 = -1.60483e-38
	(b"10000000011011110100011001011111", b"00000000000000000000000000000000"),
	(b"00000000011001110011001101010110", b"10000000000010000001001100001001"), -- -1.0219e-38 + 9.47747e-39 = -7.41512e-40
	(b"00000000011000000000011001101011", b"00000000000000000000000000000000"),
	(b"00000000000110001011000110101100", b"00000000011110001011100000010111"), -- 8.81851e-39 + 2.26779e-39 = 1.10863e-38
	(b"00000000000000100100011111001110", b"00000000000000000000000000000000"),
	(b"00000000011101010001000111111010", b"00000000011101110101100111001000"), -- 2.0943e-40 + 1.07512e-38 = 1.09606e-38
	(b"10000000000011111010100010100111", b"00000000000000000000000000000000"),
	(b"10000000011101101111101100100011", b"10000000100001101010001111001010"), -- -1.43803e-39 + -1.09267e-38 = -1.23647e-38
	(b"10000000001011000111000000000001", b"00000000000000000000000000000000"),
	(b"00000000011110000011010100011110", b"00000000010010111100010100011101"), -- -4.08094e-39 + 1.10393e-38 = 6.95837e-39
	(b"10000000001011100111010001010011", b"00000000000000000000000000000000"),
	(b"10000000001011001010001000110110", b"10000000010110110001011010001001"), -- -4.26616e-39 + -4.09895e-39 = -8.36511e-39
	(b"10000000001101111011101110101111", b"00000000000000000000000000000000"),
	(b"10000000010101111011110101000001", b"10000000100011110111100011110000"), -- -5.11828e-39 + -8.05758e-39 = -1.31759e-38
	(b"10000000010110111000100001100011", b"00000000000000000000000000000000"),
	(b"10000000011110010110101010101110", b"10000000110101001111001100010001"), -- -8.40596e-39 + -1.11504e-38 = -1.95563e-38
	(b"10000000011000001101110101110001", b"00000000000000000000000000000000"),
	(b"10000000011011110000111101111000", b"10000000110011111110110011101001"), -- -8.89565e-39 + -1.01993e-38 = -1.90949e-38
	(b"10000000001011011110111111010110", b"00000000000000000000000000000000"),
	(b"10000000000010101110111100000001", b"10000000001110001101111011010111"), -- -4.21863e-39 + -1.00409e-39 = -5.22273e-39
	(b"00000000001000111101001110000110", b"00000000000000000000000000000000"),
	(b"10000000011101000001000001101110", b"10000000010100000011110011101000"), -- 3.29012e-39 + -1.06588e-38 = -7.36869e-39
	(b"10000000000101000001011110011000", b"00000000000000000000000000000000"),
	(b"10000000011111001001011010111110", b"10000000100100001010111001010110"), -- -1.84517e-39 + -1.14417e-38 = -1.32869e-38
	(b"00000000000111101000010111010011", b"00000000000000000000000000000000"),
	(b"10000000001110110001010110111100", b"10000000000111001000111111101001"), -- 2.80307e-39 + -5.42609e-39 = -2.62302e-39
	(b"00000000011010010011100011011000", b"00000000000000000000000000000000"),
	(b"00000000000010010101010010001111", b"00000000011100101000110101100111"), -- 9.66312e-39 + 8.56853e-40 = 1.052e-38
	(b"10000000010100100111101110000010", b"00000000000000000000000000000000"),
	(b"10000000000011000101010110001100", b"10000000010111101101000100001110"), -- -7.57482e-39 + -1.13271e-39 = -8.70753e-39
	(b"00000000000111110111101101010011", b"00000000000000000000000000000000"),
	(b"10000000010000011110010001110010", b"10000000001000100110100100011111"), -- 2.89114e-39 + -6.05126e-39 = -3.16012e-39
	(b"10000000011101100111110110011011", b"00000000000000000000000000000000"),
	(b"00000000010000100010101111011001", b"10000000001101000101000111000010"), -- -1.08816e-38 + 6.07687e-39 = -4.80477e-39
	(b"00000000010001110000010101111001", b"00000000000000000000000000000000"),
	(b"10000000000010111011010110111110", b"00000000001110110100111110111011"), -- 6.52228e-39 + -1.07539e-39 = 5.4469e-39
	(b"10000000001110110111100000111001", b"00000000000000000000000000000000"),
	(b"00000000000001100101111000110110", b"10000000001101010001101000000011"), -- -5.46142e-39 + 5.84809e-40 = -4.87661e-39
	(b"00000000000001010000011000010001", b"00000000000000000000000000000000"),
	(b"00000000011010000110100000101010", b"00000000011011010110111000111011"), -- 4.61354e-40 + 9.58826e-39 = 1.00496e-38
	(b"00000000011010100100100000110100", b"00000000000000000000000000000000"),
	(b"00000000000101001100010001010011", b"00000000011111110000110010000111"), -- 9.76046e-39 + 1.90714e-39 = 1.16676e-38
	(b"10000000000100000000001000010100", b"00000000000000000000000000000000"),
	(b"10000000001000101101001101110110", b"10000000001100101101010110001010"), -- -1.47011e-39 + -3.19826e-39 = -4.66838e-39
	(b"00000000011110110001010111101100", b"00000000000000000000000000000000"),
	(b"10000000010000111011111100100110", b"00000000001101110101011011000110"), -- 1.13036e-38 + -6.22155e-39 = 5.08208e-39
	(b"00000000000000000100001011011010", b"00000000000000000000000000000000"),
	(b"10000000011100111100000000011000", b"10000000011100110111110100111110"), -- 2.39818e-41 + -1.063e-38 = -1.0606e-38
	(b"10000000000110111001110000000000", b"00000000000000000000000000000000"),
	(b"10000000011001010110101110000101", b"10000000100000010000011110000101"), -- -2.53552e-39 + -9.31396e-39 = -1.18495e-38
	(b"00000000010000101010001111011100", b"00000000000000000000000000000000"),
	(b"10000000011001011100100000110010", b"10000000001000110010010001010110"), -- 6.11992e-39 + -9.3472e-39 = -3.22728e-39
	(b"00000000001000011100110101100111", b"00000000000000000000000000000000"),
	(b"00000000010110100111110110110011", b"00000000011111000100101100011010"), -- 3.10426e-39 + 8.31029e-39 = 1.14145e-38
	(b"10000000001011010101101111100011", b"00000000000000000000000000000000"),
	(b"10000000001111001001100010111100", b"10000000011010011111010010011111"), -- -4.16556e-39 + -5.56492e-39 = -9.73048e-39
	(b"00000000010001011101000111111100", b"00000000000000000000000000000000"),
	(b"10000000000010001100101000001010", b"00000000001111010000011111110010"), -- 6.41198e-39 + -8.07162e-40 = 5.60482e-39
	(b"10000000010000100101011010001001", b"00000000000000000000000000000000"),
	(b"10000000001011100000010111110111", b"10000000011100000101110010000000"), -- -6.09219e-39 + -4.22657e-39 = -1.03188e-38
	(b"00000000001010101011101101101111", b"00000000000000000000000000000000"),
	(b"00000000001011010011110001101011", b"00000000010101111111011111011010"), -- 3.92433e-39 + 4.15427e-39 = 8.0786e-39
	(b"00000000011010011100011010111100", b"00000000000000000000000000000000"),
	(b"10000000000110110101001101110000", b"00000000010011100111001101001100"), -- 9.71402e-39 + -2.50949e-39 = 7.20453e-39
	(b"10000000010100110000100100110011", b"00000000000000000000000000000000"),
	(b"10000000000000010110010100010000", b"10000000010101000110111001000011"), -- -7.62565e-39 + -1.2809e-40 = -7.75374e-39
	(b"00000000000011011010101000101111", b"00000000000000000000000000000000"),
	(b"00000000010101011011100011010000", b"00000000011000110110001011111111"), -- 1.25491e-39 + 7.87232e-39 = 9.12723e-39
	(b"00000000011111000000001110110000", b"00000000000000000000000000000000"),
	(b"00000000010001010011011011001111", b"00000000110000010011101001111111"), -- 1.13889e-38 + 6.35631e-39 = 1.77452e-38
	(b"10000000000101011010011100011111", b"00000000000000000000000000000000"),
	(b"10000000001000011010100001100110", b"10000000001101110100111110000101"), -- -1.9885e-39 + -3.09098e-39 = -5.07948e-39
	(b"00000000011101100011100010101000", b"00000000000000000000000000000000"),
	(b"10000000001000000000100001111100", b"00000000010101100011000000101100"), -- 1.08569e-38 + -2.94178e-39 = 7.91513e-39
	(b"10000000011001100110100010000100", b"00000000000000000000000000000000"),
	(b"10000000011001010110110110100011", b"10000000110010111101011000100111"), -- -9.40471e-39 + -9.31472e-39 = -1.87194e-38
	(b"00000000000100100001011001000110", b"00000000000000000000000000000000"),
	(b"10000000000100111000010010100110", b"10000000000000010110111001100000"), -- 1.66103e-39 + -1.79246e-39 = -1.31431e-40
	(b"10000000010111101101000000010100", b"00000000000000000000000000000000"),
	(b"00000000010111101111101110011111", b"00000000000000000010101110001011"), -- -8.70718e-39 + 8.7228e-39 = 1.56203e-41
	(b"10000000000100101100000001000101", b"00000000000000000000000000000000"),
	(b"10000000011101101100000110110110", b"10000000100010011000000111111011"), -- -1.72201e-39 + -1.09061e-38 = -1.26281e-38
	(b"10000000011111000011100100100111", b"00000000000000000000000000000000"),
	(b"10000000000101001010100000101001", b"10000000100100001110000101010000"), -- -1.14081e-38 + -1.89703e-39 = -1.33051e-38
	(b"00000000001111000001010000000000", b"00000000000000000000000000000000"),
	(b"00000000010100111010001111110011", b"00000000100011111011011111110011"), -- 5.5173e-39 + 7.68116e-39 = 1.31985e-38
	(b"00000000010001010111000101110110", b"00000000000000000000000000000000"),
	(b"10000000011101011101101010000011", b"10000000001100000110100100001101"), -- 6.37735e-39 + -1.08231e-38 = -4.44579e-39
	(b"00000000001010010010101111010100", b"00000000000000000000000000000000"),
	(b"00000000011001100111011010010001", b"00000000100011111010001001100101"), -- 3.78098e-39 + 9.40975e-39 = 1.31907e-38
	(b"10000000001101101101000000001100", b"00000000000000000000000000000000"),
	(b"10000000011111010110111101111011", b"10000000101101000011111110000111"), -- -5.03375e-39 + -1.15194e-38 = -1.65532e-38
	(b"10000000001011110110000100100101", b"00000000000000000000000000000000"),
	(b"00000000011010000110011100100000", b"00000000001110010000010111111011"), -- -4.35112e-39 + 9.58789e-39 = 5.23677e-39
	(b"10000000000110010000111101001010", b"00000000000000000000000000000000"),
	(b"00000000011010111101100111011011", b"00000000010100101100101010010001"), -- -2.30137e-39 + 9.90455e-39 = 7.60318e-39
	(b"10000000010001010010100110111100", b"00000000000000000000000000000000"),
	(b"10000000000011010100000011001101", b"10000000010100100110101010001001"), -- -6.35162e-39 + -1.21711e-39 = -7.56873e-39
	(b"10000000001000000100001111011011", b"00000000000000000000000000000000"),
	(b"00000000011101111000011010101001", b"00000000010101110100001011001110"), -- -2.96308e-39 + 1.09767e-38 = 8.01365e-39
	(b"10000000011010111010000111101011", b"00000000000000000000000000000000"),
	(b"10000000011011000100101011101010", b"10000000110101111110110011010101"), -- -9.88448e-39 + -9.94511e-39 = -1.98296e-38
	(b"00000000001000010001111000111001", b"00000000000000000000000000000000"),
	(b"10000000010101000100111001000000", b"10000000001100110011000000000111"), -- 3.04141e-39 + -7.74225e-39 = -4.70084e-39
	(b"00000000000001001011000010000010", b"00000000000000000000000000000000"),
	(b"00000000000001000011111001001011", b"00000000000010001110111011001101"), -- 4.30661e-40 + 3.89688e-40 = 8.2035e-40
	(b"00000000000110110011100110000110", b"00000000000000000000000000000000"),
	(b"10000000001100101011111011010101", b"10000000000101111000010101001111"), -- 2.50019e-39 + -4.66023e-39 = -2.16004e-39
	(b"00000000001011010010101011011100", b"00000000000000000000000000000000"),
	(b"10000000000011101010010110100100", b"00000000000111101000010100111000"), -- 4.14797e-39 + -1.34512e-39 = 2.80285e-39
	(b"00000000011001101100010011110011", b"00000000000000000000000000000000"),
	(b"10000000011111000110011100001110", b"10000000000101011010001000011011"), -- 9.43787e-39 + -1.14246e-38 = -1.9867e-39
	(b"00000000010111011001101010001110", b"00000000000000000000000000000000"),
	(b"00000000001010011111111010101110", b"00000000100001111001100100111100"), -- 8.59614e-39 + 3.85662e-39 = 1.24528e-38
	(b"00000000011111100010001110111000", b"00000000000000000000000000000000"),
	(b"10000000010000111110000000101100", b"00000000001110100100001110001100"), -- 1.15841e-38 + -6.2334e-39 = 5.35069e-39
	(b"10000000011010111101010000111011", b"00000000000000000000000000000000"),
	(b"10000000000110101011001011100011", b"10000000100001101000011100011110"), -- -9.90253e-39 + -2.4519e-39 = -1.23544e-38
	(b"10000000011101111110000111100110", b"00000000000000000000000000000000"),
	(b"10000000010101010111110110110101", b"10000000110011010101111110011011"), -- -1.10095e-38 + -7.85111e-39 = -1.88606e-38
	(b"10000000001011000110001011100101", b"00000000000000000000000000000000"),
	(b"10000000010111000100100000111000", b"10000000100010001010101100011101"), -- -4.07624e-39 + -8.47477e-39 = -1.2551e-38
	(b"00000000011000110000000001101111", b"00000000000000000000000000000000"),
	(b"10000000011110111111000001110011", b"10000000000110001111000000000100"), -- 9.09187e-39 + -1.1382e-38 = -2.29015e-39
	(b"00000000010011111000111100100001", b"00000000000000000000000000000000"),
	(b"00000000010011101000001011100111", b"00000000100111100001001000001000"), -- 7.30635e-39 + 7.21013e-39 = 1.45165e-38
	(b"00000000011000010101001110100000", b"00000000000000000000000000000000"),
	(b"00000000011011010001011111010110", b"00000000110011100110101101110110"), -- 8.93804e-39 + 1.00186e-38 = 1.89567e-38
	(b"10000000001010101101100111010101", b"00000000000000000000000000000000"),
	(b"10000000000110010000111011001101", b"10000000010000111110100010100010"), -- -3.93523e-39 + -2.3012e-39 = -6.23643e-39
	(b"00000000000001000110000100001100", b"00000000000000000000000000000000"),
	(b"00000000000011101011110000110011", b"00000000000100110001110100111111"), -- 4.02156e-40 + 1.35321e-39 = 1.75537e-39
	(b"00000000000110001000101110001101", b"00000000000000000000000000000000"),
	(b"10000000001110000111011011000000", b"10000000000111111110101100110011"), -- 2.25411e-39 + -5.18539e-39 = -2.93127e-39
	(b"10000000010100010000110010111010", b"00000000000000000000000000000000"),
	(b"10000000000000001110101100000010", b"10000000010100011111011110111100"), -- -7.44324e-39 + -8.43049e-41 = -7.52755e-39
	(b"10000000010100011101110111000000", b"00000000000000000000000000000000"),
	(b"00000000001001010010010010100111", b"10000000001011001011100100011001"), -- -7.51822e-39 + 3.41106e-39 = -4.10716e-39
	(b"10000000011101001011001011010101", b"00000000000000000000000000000000"),
	(b"10000000010100110001110001111011", b"10000000110001111100111101010000"), -- -1.07171e-38 + -7.63256e-39 = -1.83496e-38
	(b"00000000011101101111001111110110", b"00000000000000000000000000000000"),
	(b"10000000010010100000100110100101", b"00000000001011001110101001010001"), -- 1.09241e-38 + -6.79929e-39 = 4.12482e-39
	(b"00000000011000101111001010100101", b"00000000000000000000000000000000"),
	(b"10000000001101000110000011111011", b"00000000001011101001000110101010"), -- 9.08692e-39 + -4.81024e-39 = 4.27669e-39
	(b"00000000010001011000000101010101", b"00000000000000000000000000000000"),
	(b"10000000001110011110110111000000", b"00000000000010111001001110010101"), -- 6.38304e-39 + -5.31991e-39 = 1.06313e-39
	(b"10000000010010110001001100011010", b"00000000000000000000000000000000"),
	(b"00000000000101010001001010011000", b"10000000001101100000000010000010"), -- -6.89451e-39 + 1.93522e-39 = -4.9593e-39
	(b"00000000011100111101110010010110", b"00000000000000000000000000000000"),
	(b"00000000001001100000101101111101", b"00000000100110011110100000010011"), -- 1.06402e-38 + 3.49387e-39 = 1.41341e-38
	(b"10000000010001011100110110100110", b"00000000000000000000000000000000"),
	(b"00000000000011110011101101010001", b"10000000001101101001001001010101"), -- -6.41042e-39 + 1.39881e-39 = -5.01161e-39
	(b"00000000010101101110000111101111", b"00000000000000000000000000000000"),
	(b"00000000001110110001111101100101", b"00000000100100100000000101010100"), -- 7.9789e-39 + 5.42956e-39 = 1.34085e-38
	(b"00000000011110111001110111110111", b"00000000000000000000000000000000"),
	(b"00000000011110101110001010010101", b"00000000111101101000000010001100"), -- 1.13524e-38 + 1.12852e-38 = 2.26376e-38
	(b"00000000001101101000111101100101", b"00000000000000000000000000000000"),
	(b"00000000011010110011011010110111", b"00000000101000011100011000011100"), -- 5.01056e-39 + 9.84603e-39 = 1.48566e-38
	(b"00000000010100111110101100100001", b"00000000000000000000000000000000"),
	(b"00000000010000001010100000111110", b"00000000100101001001001101011111"), -- 7.70669e-39 + 5.93783e-39 = 1.36445e-38
	(b"00000000010010110101011111110100", b"00000000000000000000000000000000"),
	(b"10000000011001100110100010101100", b"10000000000110110001000010111000"), -- 6.91921e-39 + -9.40477e-39 = -2.48556e-39
	(b"00000000010100001100101110111110", b"00000000000000000000000000000000"),
	(b"10000000010110010100111100010010", b"10000000000010001000001101010100"), -- 7.41993e-39 + -8.20172e-39 = -7.81796e-40
	(b"00000000010100010011100111101111", b"00000000000000000000000000000000"),
	(b"00000000010101000101010000110010", b"00000000101001011000111000100001"), -- 7.45946e-39 + 7.74439e-39 = 1.52038e-38
	(b"10000000011111100110110001111000", b"00000000000000000000000000000000"),
	(b"00000000001010101111011010011011", b"10000000010100110111010111011101"), -- -1.16102e-38 + 3.94556e-39 = -7.66463e-39
	(b"10000000011000011100010101010000", b"00000000000000000000000000000000"),
	(b"00000000011111110001001101000110", b"00000000000111010100110111110110"), -- -8.97883e-39 + 1.167e-38 = 2.6912e-39
	(b"10000000010010000001100011010111", b"00000000000000000000000000000000"),
	(b"10000000011011100010101000001001", b"10000000101101100100001011100000"), -- -6.62107e-39 + -1.0117e-38 = -1.67381e-38
	(b"10000000011001110101101101011010", b"00000000000000000000000000000000"),
	(b"10000000001111111100101010010011", b"10000000101001110010010111101101"), -- -9.49183e-39 + -5.85831e-39 = -1.53501e-38
	(b"00000000010001110100100110010110", b"00000000000000000000000000000000"),
	(b"10000000000101011011000010100110", b"00000000001100011001100011110000"), -- 6.54672e-39 + -1.99191e-39 = 4.5548e-39
	(b"10000000011010100011110100110111", b"00000000000000000000000000000000"),
	(b"00000000011100101000100100111100", b"00000000000010000100110000000101"), -- -9.75652e-39 + 1.05185e-38 = 7.61955e-40
	(b"10000000010101001111011100111100", b"00000000000000000000000000000000"),
	(b"00000000000110011001101111000000", b"10000000001110110101101101111100"), -- -7.80287e-39 + 2.35176e-39 = -5.45111e-39
	(b"00000000010010011000011010101111", b"00000000000000000000000000000000"),
	(b"00000000011110011001110001010110", b"00000000110000110010001100000101"), -- 6.75231e-39 + 1.11682e-38 = 1.79205e-38
	(b"10000000000100010000010001110010", b"00000000000000000000000000000000"),
	(b"00000000001001010000010011110011", b"00000000000101000000000010000001"), -- -1.5628e-39 + 3.39969e-39 = 1.83689e-39
	(b"00000000001100001010110000010001", b"00000000000000000000000000000000"),
	(b"00000000011010100000111011011111", b"00000000100110101011101011110000"), -- 4.46983e-39 + 9.7399e-39 = 1.42097e-38
	(b"00000000001111011110111000110000", b"00000000000000000000000000000000"),
	(b"00000000000000001111010101111111", b"00000000001111101110001110101111"), -- 5.68741e-39 + 8.80674e-41 = 5.77548e-39
	(b"10000000000101100010110110010111", b"00000000000000000000000000000000"),
	(b"10000000011111110011000001110010", b"10000000100101010101111000001001"), -- -2.03674e-39 + -1.16805e-38 = -1.37172e-38
	(b"00000000000000011111001101100110", b"00000000000000000000000000000000"),
	(b"10000000010100111101101101111000", b"10000000010100011110100000010010"), -- 1.7915e-40 + -7.70108e-39 = -7.52193e-39
	(b"00000000011011001111010100101100", b"00000000000000000000000000000000"),
	(b"00000000001101110010000000101110", b"00000000101001000001010101011010"), -- 1.00062e-38 + 5.0625e-39 = 1.50687e-38
	(b"10000000001101100001100100000101", b"00000000000000000000000000000000"),
	(b"10000000000100110010001100100001", b"10000000010010010011110000100110"), -- -4.96809e-39 + -1.75748e-39 = -6.72557e-39
	(b"10000000010110110101001100100011", b"00000000000000000000000000000000"),
	(b"00000000000000001110100110101011", b"10000000010110100110100101111000"), -- -8.38685e-39 + 8.38243e-41 = -8.30303e-39
	(b"10000000010001101001001001111011", b"00000000000000000000000000000000"),
	(b"10000000001011101101101100111011", b"10000000011101010110110110110110"), -- -6.48103e-39 + -4.30308e-39 = -1.07841e-38
	(b"10000000011110111000001000110010", b"00000000000000000000000000000000"),
	(b"10000000000111111110111011110000", b"10000000100110110111000100100010"), -- -1.13425e-38 + -2.93262e-39 = -1.42751e-38
	(b"10000000001001111101111100000000", b"00000000000000000000000000000000"),
	(b"10000000011100110000011110010101", b"10000000100110101110011010010101"), -- -3.66158e-39 + -1.05638e-38 = -1.42254e-38
	(b"10000000010010110010010100110010", b"00000000000000000000000000000000"),
	(b"10000000000100101001110010000100", b"10000000010111011100000110110110"), -- -6.90101e-39 + -1.70919e-39 = -8.61019e-39
	(b"10000000000111011100010100000011", b"00000000000000000000000000000000"),
	(b"10000000001111011101011110100111", b"10000000010110111001110010101010"), -- -2.7339e-39 + -5.67933e-39 = -8.41323e-39
	(b"10000000011101101100100101011011", b"00000000000000000000000000000000"),
	(b"10000000000000111011011010111101", b"10000000011110101000000000011000"), -- -1.09088e-38 + -3.41061e-40 = -1.12499e-38
	(b"10000000001000000000110010010100", b"00000000000000000000000000000000"),
	(b"00000000011100000101000100000101", b"00000000010100000100010001110001"), -- -2.94325e-39 + 1.03146e-38 = 7.37139e-39
	(b"10000000000110100001001010011000", b"00000000000000000000000000000000"),
	(b"10000000001001001011101111100101", b"10000000001111101100111001111101"), -- -2.39439e-39 + -3.37348e-39 = -5.76787e-39
	(b"10000000010001000111011111011101", b"00000000000000000000000000000000"),
	(b"00000000011010011011011000010001", b"00000000001001010011111000110100"), -- -6.28781e-39 + 9.70804e-39 = 3.42023e-39
	(b"00000000000101001101110010101100", b"00000000000000000000000000000000"),
	(b"00000000011000010001101000111000", b"00000000011101011111011011100100"), -- 1.91587e-39 + 8.91745e-39 = 1.08333e-38
	(b"00000000001111001100000011000011", b"00000000000000000000000000000000"),
	(b"10000000001110100111111011000000", b"00000000000000100100001000000011"), -- 5.57928e-39 + -5.37193e-39 = 2.07352e-40
	(b"00000000011100010100101101111000", b"00000000000000000000000000000000"),
	(b"10000000011111100001001001000100", b"10000000000011001100011011001100"), -- 1.04045e-38 + -1.15778e-38 = -1.17334e-39
	(b"10000000010010001001111110100001", b"00000000000000000000000000000000"),
	(b"10000000000111011100010011110001", b"10000000011001100110010010010010"), -- -6.66942e-39 + -2.73388e-39 = -9.4033e-39
	(b"00000000001111110100101000011011", b"00000000000000000000000000000000"),
	(b"00000000000011110100011010000001", b"00000000010011101001000010011100"), -- 5.81222e-39 + 1.40282e-39 = 7.21504e-39
	(b"00000000000011101110011010010001", b"00000000000000000000000000000000"),
	(b"00000000010100011011101001100010", b"00000000011000001010000011110011"), -- 1.36841e-39 + 7.50554e-39 = 8.87395e-39
	(b"10000000000101001000101001110000", b"00000000000000000000000000000000"),
	(b"10000000000001000111100110101100", b"10000000000110010000010000011100"), -- -1.88637e-39 + -4.1099e-40 = -2.29736e-39
	(b"00000000000100010101011101010010", b"00000000000000000000000000000000"),
	(b"00000000000101100000111001011001", b"00000000001001110110010110101011"), -- 1.59253e-39 + 2.02553e-39 = 3.61806e-39
	(b"00000000000000010001010010011110", b"00000000000000000000000000000000"),
	(b"10000000010100010111001001000011", b"10000000010100000101110110100101"), -- 9.92315e-41 + -7.47966e-39 = -7.38043e-39
	(b"00000000001001110010111010111101", b"00000000000000000000000000000000"),
	(b"10000000001111000001000000010001", b"10000000000101001110000101010100"), -- 3.59835e-39 + -5.51589e-39 = -1.91754e-39
	(b"10000000011101100100110100101011", b"00000000000000000000000000000000"),
	(b"10000000011111111000011100010100", b"10000000111101011101010000111111"), -- -1.08643e-38 + -1.17116e-38 = -2.25758e-38
	(b"10000000011110000111100011001010", b"00000000000000000000000000000000"),
	(b"10000000010101011100001111100001", b"10000000110011100011110010101011"), -- -1.10636e-38 + -7.87629e-39 = -1.89399e-38
	(b"00000000000110100100100010111001", b"00000000000000000000000000000000"),
	(b"10000000001000000111111100000110", b"10000000000001100011011001001101"), -- 2.41381e-39 + -2.9843e-39 = -5.70492e-40
	(b"10000000000001011011010011011101", b"00000000000000000000000000000000"),
	(b"10000000010101101100111111111100", b"10000000010111001000010011011001"), -- -5.24059e-40 + -7.97246e-39 = -8.49652e-39
	(b"10000000010001000100110111011111", b"00000000000000000000000000000000"),
	(b"10000000000101101110101010000101", b"10000000010110110011100001100100"), -- -6.27275e-39 + -2.10451e-39 = -8.37726e-39
	(b"10000000010110111001001001000011", b"00000000000000000000000000000000"),
	(b"10000000001010010010111010100000", b"10000000100001001100000011100011"), -- -8.4095e-39 + -3.78198e-39 = -1.21915e-38
	(b"10000000011000000001110100101101", b"00000000000000000000000000000000"),
	(b"10000000000111010001111101001001", b"10000000011111010011110001110110"), -- -8.82667e-39 + -2.67445e-39 = -1.15011e-38
	(b"00000000011100111001111011010010", b"00000000000000000000000000000000"),
	(b"00000000000000110010101000001011", b"00000000011101101100100011011101"), -- 1.06181e-38 + 2.90589e-40 = 1.09086e-38
	(b"00000000010000100100000101010001", b"00000000000000000000000000000000"),
	(b"10000000001000011100011111111010", b"00000000001000000111100101010111"), -- 6.08457e-39 + -3.10231e-39 = 2.98226e-39
	(b"00000000001010100000011001110110", b"00000000000000000000000000000000"),
	(b"10000000011000110110100011100010", b"10000000001110010110001001101100"), -- 3.85941e-39 + -9.12934e-39 = -5.26993e-39
	(b"10000000011000010010110001011011", b"00000000000000000000000000000000"),
	(b"00000000010001000100011101000000", b"10000000000111001110010100011011"), -- -8.92395e-39 + 6.27037e-39 = -2.65358e-39
	(b"00000000001100000100111100000101", b"00000000000000000000000000000000"),
	(b"10000000001100101101010001111101", b"10000000000000101000010101111000"), -- 4.43645e-39 + -4.668e-39 = -2.31551e-40
	(b"00000000000010111001010000011001", b"00000000000000000000000000000000"),
	(b"10000000010110100101011110100000", b"10000000010011101100001110000111"), -- 1.06332e-39 + -8.29663e-39 = -7.23331e-39
	(b"00000000001001101101111000100111", b"00000000000000000000000000000000"),
	(b"00000000011001101100000001011101", b"00000000100011011001111010000100"), -- 3.56944e-39 + 9.43623e-39 = 1.30057e-38
	(b"10000000010011010111001001101010", b"00000000000000000000000000000000"),
	(b"10000000000010110111000010111010", b"10000000010110001110001100100100"), -- -7.11238e-39 + -1.05063e-39 = -8.16301e-39
	(b"10000000010011011010101000110001", b"00000000000000000000000000000000"),
	(b"00000000011111111111001110011001", b"00000000001100100100100101101000"), -- -7.13239e-39 + 1.17505e-38 = 4.61811e-39
	(b"10000000011010101100110100010111", b"00000000000000000000000000000000"),
	(b"10000000000100101001010101001110", b"10000000011111010110001001100101"), -- -9.80813e-39 + -1.7066e-39 = -1.15147e-38
	(b"10000000001111001000100101000011", b"00000000000000000000000000000000"),
	(b"00000000011001110101000111110101", b"00000000001010101100100010110010"), -- -5.55937e-39 + 9.48846e-39 = 3.92909e-39
	(b"10000000011101111111100010000111", b"00000000000000000000000000000000"),
	(b"10000000010111001101011101110010", b"10000000110101001100111111111001"), -- -1.10176e-38 + -8.52615e-39 = -1.95437e-38
	(b"00000000011001010110000100111001", b"00000000000000000000000000000000"),
	(b"00000000000111110000101011001101", b"00000000100001000110110000000110"), -- 9.31026e-39 + 2.85077e-39 = 1.2161e-38
	(b"00000000011001011100010110011001", b"00000000000000000000000000000000"),
	(b"10000000011101111101110001010001", b"10000000000100100001011010111000"), -- 9.34627e-39 + -1.10075e-38 = -1.66119e-39
	(b"10000000010101001101111101000110", b"00000000000000000000000000000000"),
	(b"00000000010110000000011010111010", b"00000000000000110010011101110100"), -- -7.79428e-39 + 8.08394e-39 = 2.8966e-40
	(b"10000000000001111100101001111011", b"00000000000000000000000000000000"),
	(b"00000000010001011111101000011111", b"00000000001111100010111110100100"), -- -7.15485e-40 + 6.42638e-39 = 5.71089e-39
	(b"10000000001010101001100011000000", b"00000000000000000000000000000000"),
	(b"10000000001110111111001011101001", b"10000000011001101000101110101001"), -- -3.91189e-39 + -5.50543e-39 = -9.41732e-39
	(b"00000000010001000000000101111010", b"00000000000000000000000000000000"),
	(b"00000000010101110011101101100101", b"00000000100110110011110011011111"), -- 6.24534e-39 + 8.01099e-39 = 1.42563e-38
	(b"10000000001001110010000001000001", b"00000000000000000000000000000000"),
	(b"10000000011011011110011101110001", b"10000000100101010000011110110010"), -- -3.59315e-39 + -1.00931e-38 = -1.36862e-38
	(b"00000000000011000000011001000000", b"00000000000000000000000000000000"),
	(b"10000000001000010110111100011100", b"10000000000101010110100011011100"), -- 1.10427e-39 + -3.07043e-39 = -1.96616e-39
	(b"00000000011100101100110001001011", b"00000000000000000000000000000000"),
	(b"00000000011001110010001111111110", b"00000000110110011111000001001001"), -- 1.05425e-38 + 9.47197e-39 = 2.00145e-38
	(b"00000000001010010100001110100111", b"00000000000000000000000000000000"),
	(b"10000000010001111001010101000100", b"10000000000111100101000110011101"), -- 3.78952e-39 + -6.57387e-39 = -2.78434e-39
	(b"00000000001110001101111111000000", b"00000000000000000000000000000000"),
	(b"00000000010111001001111001010010", b"00000000100101010111111000010010"), -- 5.22305e-39 + 8.50566e-39 = 1.37287e-38
	(b"00000000000100111011110101101011", b"00000000000000000000000000000000"),
	(b"10000000010011000100110001101111", b"10000000001110001000111100000100"), -- 1.81282e-39 + -7.00692e-39 = -5.19409e-39
	(b"00000000000110011110000011011100", b"00000000000000000000000000000000"),
	(b"00000000011001111001000101000100", b"00000000100000010111001000100000"), -- 2.37655e-39 + 9.51117e-39 = 1.18877e-38
	(b"10000000001101110101000110000001", b"00000000000000000000000000000000"),
	(b"10000000010101100111101110110110", b"10000000100011011100110100110111"), -- -5.08019e-39 + -7.94223e-39 = -1.30224e-38
	(b"10000000010100110011000001011101", b"00000000000000000000000000000000"),
	(b"10000000010011000111111001010110", b"10000000100111111010111010110011"), -- -7.6397e-39 + -7.02482e-39 = -1.46645e-38
	(b"00000000011100010110000110000101", b"00000000000000000000000000000000"),
	(b"00000000000011001100000101011101", b"00000000011111100010001011100010"), -- 1.04124e-38 + 1.17139e-39 = 1.15838e-38
	(b"00000000000001000111001001100001", b"00000000000000000000000000000000"),
	(b"00000000001010001100101010100010", b"00000000001011010011110100000011"), -- 4.08373e-40 + 3.74611e-39 = 4.15448e-39
	(b"00000000000010111000101100100011", b"00000000000000000000000000000000"),
	(b"00000000000000111101001101011000", b"00000000000011110101111001111011"), -- 1.0601e-39 + 3.51322e-40 = 1.41143e-39
	(b"00000000011101000001110110000101", b"00000000000000000000000000000000"),
	(b"10000000010001101111100110111100", b"00000000001011010010001111001001"), -- 1.06635e-38 + -6.51807e-39 = 4.14543e-39
	(b"10000000010100001110110110111110", b"00000000000000000000000000000000"),
	(b"00000000011111010111110011011100", b"00000000001011001000111100011110"), -- -7.43213e-39 + 1.15242e-38 = 4.0921e-39
	(b"00000000011000001001010101110101", b"00000000000000000000000000000000"),
	(b"00000000000010110110101011000000", b"00000000011011000000000000110101"), -- 8.86982e-39 + 1.04849e-39 = 9.91831e-39
	(b"10000000011001111110011000011110", b"00000000000000000000000000000000"),
	(b"00000000000000100101000011011010", b"10000000011001011001010101000100"), -- -9.54161e-39 + 2.12675e-40 = -9.32893e-39
	(b"10000000010000001010100011101001", b"00000000000000000000000000000000"),
	(b"10000000011111001001110100011011", b"10000000101111010100011000000100"), -- -5.93807e-39 + -1.1444e-38 = -1.7382e-38
	(b"10000000001010110110010001110011", b"00000000000000000000000000000000"),
	(b"10000000001110010010110011100001", b"10000000011001001001000101010100"), -- -3.98496e-39 + -5.25072e-39 = -9.23568e-39
	(b"10000000010010010101010110011000", b"00000000000000000000000000000000"),
	(b"10000000001100101001001110101000", b"10000000011110111110100101000000"), -- -6.7347e-39 + -4.64474e-39 = -1.13794e-38
	(b"10000000001111001011010001011110", b"00000000000000000000000000000000"),
	(b"10000000001100011101110001001001", b"10000000011011101001000010100111"), -- -5.57483e-39 + -4.57896e-39 = -1.01538e-38
	(b"10000000010100100011111010000000", b"00000000000000000000000000000000"),
	(b"00000000011011111111110111010000", b"00000000000111011011111101010000"), -- -7.55293e-39 + 1.02848e-38 = 2.73186e-39
	(b"10000000000100000110111100010011", b"00000000000000000000000000000000"),
	(b"00000000011111011001010100000100", b"00000000011011010010010111110001"), -- -1.50921e-39 + 1.15329e-38 = 1.00237e-38
	(b"00000000001111111111010110100000", b"00000000000000000000000000000000"),
	(b"00000000001111000000001100100101", b"00000000011110111111100011000101"), -- 5.87375e-39 + 5.51126e-39 = 1.1385e-38
	(b"00000000010101110010111010001100", b"00000000000000000000000000000000"),
	(b"00000000010100010000001000000001", b"00000000101010000011000010001101"), -- 8.00639e-39 + 7.43939e-39 = 1.54458e-38
	(b"00000000001110000100011011011110", b"00000000000000000000000000000000"),
	(b"00000000010101100111110101010010", b"00000000100011101100010000110000"), -- 5.16821e-39 + 7.94281e-39 = 1.3111e-38
	(b"10000000000100000000101100111111", b"00000000000000000000000000000000"),
	(b"00000000011001011001011011011111", b"00000000010101011000101110100000"), -- -1.4734e-39 + 9.32951e-39 = 7.85611e-39
	(b"10000000010001101110001111001000", b"00000000000000000000000000000000"),
	(b"10000000011000001001000010000000", b"10000000101001110111010001001000"), -- -6.5102e-39 + -8.86804e-39 = -1.53782e-38
	(b"10000000000110100011100100000111", b"00000000000000000000000000000000"),
	(b"10000000001010110000000101010111", b"10000000010001010011101001011110"), -- -2.40818e-39 + -3.94941e-39 = -6.35759e-39
	(b"00000000000001011011111111010011", b"00000000000000000000000000000000"),
	(b"10000000011111101111001101111001", b"10000000011110010011001110100110"), -- 5.27991e-40 + -1.16586e-38 = -1.11306e-38
	(b"00000000000000011000110111100001", b"00000000000000000000000000000000"),
	(b"00000000010001101000100011100100", b"00000000010010000001011011000101"), -- 1.42732e-40 + 6.47759e-39 = 6.62032e-39
	(b"00000000001101011101111011110110", b"00000000000000000000000000000000"),
	(b"10000000010000001110010000011001", b"10000000000010110000010100100011"), -- 4.94726e-39 + -5.9593e-39 = -1.01203e-39
	(b"10000000010101111100001001111101", b"00000000000000000000000000000000"),
	(b"10000000000010001010010001101011", b"10000000011000000110011011101000"), -- -8.05946e-39 + -7.93666e-40 = -8.85312e-39
	(b"10000000010011100001101000001101", b"00000000000000000000000000000000"),
	(b"00000000011000101111000110101110", b"00000000000101001101011110100001"), -- -7.17251e-39 + 9.08658e-39 = 1.91406e-39
	(b"00000000011000111111110010000100", b"00000000000000000000000000000000"),
	(b"10000000001010101010001111001011", b"00000000001110010101100010111001"), -- 9.1823e-39 + -3.91585e-39 = 5.26645e-39
	(b"00000000000110100110001101011010", b"00000000000000000000000000000000"),
	(b"10000000011011100011000100011101", b"10000000010100111100110111000011"), -- 2.42336e-39 + -1.01195e-38 = -7.69616e-39
	(b"10000000010010011011001010000000", b"00000000000000000000000000000000"),
	(b"00000000011100010111001101101110", b"00000000001001111100000011101110"), -- -6.76802e-39 + 1.04188e-38 = 3.65079e-39
	(b"00000000000001011010100001101111", b"00000000000000000000000000000000"),
	(b"10000000011001111010110111100010", b"10000000011000100000010101110011"), -- 5.196e-40 + -9.52143e-39 = -9.00183e-39
	(b"00000000000110000010001011001001", b"00000000000000000000000000000000"),
	(b"10000000010000110100100101100001", b"10000000001010110010011010011000"), -- 2.21653e-39 + -6.1793e-39 = -3.96277e-39
	(b"00000000011101001011011011100010", b"00000000000000000000000000000000"),
	(b"00000000000011011101000101000010", b"00000000100000101000100000100100"), -- 1.07185e-38 + 1.26893e-39 = 1.19875e-38
	(b"10000000000101011100000110111000", b"00000000000000000000000000000000"),
	(b"00000000001101100100001111010001", b"00000000001000001000001000011001"), -- -1.99804e-39 + 4.98344e-39 = 2.98541e-39
	(b"10000000011010011000011010100100", b"00000000000000000000000000000000"),
	(b"00000000010111100010001011111110", b"10000000000010110110001110100110"), -- -9.69103e-39 + 8.64509e-39 = -1.04594e-39
	(b"10000000000000101001001010001111", b"00000000000000000000000000000000"),
	(b"00000000001000101001010101101010", b"00000000001000000000001011011011"), -- -2.36246e-40 + 3.17601e-39 = 2.93976e-39
	(b"10000000000111001101110100011100", b"00000000000000000000000000000000"),
	(b"00000000011111000110000110011100", b"00000000010111111000010010000000"), -- -2.65071e-39 + 1.14226e-38 = 8.7719e-39
	(b"00000000000101010001000110110101", b"00000000000000000000000000000000"),
	(b"10000000010010110110100010011100", b"10000000001101100101011011100111"), -- 1.9349e-39 + -6.92519e-39 = -4.99029e-39
	(b"10000000000011010010011100011011", b"00000000000000000000000000000000"),
	(b"10000000011010000100001000000101", b"10000000011101010110100100100000"), -- -1.20789e-39 + -9.57457e-39 = -1.07825e-38
	(b"10000000001101111111001111010101", b"00000000000000000000000000000000"),
	(b"00000000001010111010100001110101", b"10000000000011000100101101100000"), -- -5.13842e-39 + 4.00936e-39 = -1.12907e-39
	(b"10000000000001010010011100000101", b"00000000000000000000000000000000"),
	(b"00000000001111001001010011011101", b"00000000001101110110110111011000"), -- -4.73175e-40 + 5.56353e-39 = 5.09036e-39
	(b"00000000000100111000101001100111", b"00000000000000000000000000000000"),
	(b"10000000001110000111000111000101", b"10000000001001001110011101011110"), -- 1.79452e-39 + -5.1836e-39 = -3.38908e-39
	(b"10000000001101000111000110011111", b"00000000000000000000000000000000"),
	(b"00000000001010010100001101001111", b"10000000000010110010111001010000"), -- -4.81621e-39 + 3.7894e-39 = -1.0268e-39
	(b"10000000011001100100101001111010", b"00000000000000000000000000000000"),
	(b"00000000010110111101001001100110", b"10000000000010100111100000010100"), -- -9.39394e-39 + 8.43251e-39 = -9.61431e-40
	(b"00000000011001000101001110011011", b"00000000000000000000000000000000"),
	(b"00000000001011001111011000011111", b"00000000100100010100100110111010"), -- 9.21354e-39 + 4.12905e-39 = 1.33426e-38
	(b"10000000011101110100001101110110", b"00000000000000000000000000000000"),
	(b"10000000000000101101100010010010", b"10000000011110100001110000001000"), -- -1.09526e-38 + -2.61362e-40 = -1.1214e-38
	(b"00000000000010101000011000110110", b"00000000000000000000000000000000"),
	(b"00000000000101110111000010101011", b"00000000001000011111011011100001"), -- 9.66501e-40 + 2.15263e-39 = 3.11913e-39
	(b"10000000010110100000011010000110", b"00000000000000000000000000000000"),
	(b"00000000000001010111100100001110", b"10000000010101001000110101111000"), -- -8.26753e-39 + 5.02604e-40 = -7.76493e-39
	(b"10000000011100000011111111000101", b"00000000000000000000000000000000"),
	(b"10000000011000110010100101110110", b"10000000110100110110100100111011"), -- -1.03085e-38 + -9.10659e-39 = -1.9415e-38
	(b"00000000001000010100010111011111", b"00000000000000000000000000000000"),
	(b"10000000011000010010000111101010", b"10000000001111111101110000001011"), -- 3.05564e-39 + -8.92021e-39 = -5.86457e-39
	(b"10000000001011110010110000001001", b"00000000000000000000000000000000"),
	(b"10000000000001000101010010011101", b"10000000001100111000000010100110"), -- -4.33207e-39 + -3.97696e-40 = -4.72976e-39
	(b"10000000001100010001011001111100", b"00000000000000000000000000000000"),
	(b"00000000010001101000100000010100", b"00000000000101010111000110011000"), -- -4.50801e-39 + 6.4773e-39 = 1.9693e-39
	(b"10000000011101101111101001110011", b"00000000000000000000000000000000"),
	(b"10000000001010010011100010101010", b"10000000101000000011001100011101"), -- -1.09264e-38 + -3.78558e-39 = -1.4712e-38
	(b"00000000011010010011010110001101", b"00000000000000000000000000000000"),
	(b"00000000011011110010000101000110", b"00000000110110000101011011010011"), -- 9.66194e-39 + 1.02057e-38 = 1.98676e-38
	(b"10000000000111000110110011111010", b"00000000000000000000000000000000"),
	(b"10000000010000101101101001011100", b"10000000010111110100011101010110"), -- -2.61049e-39 + -6.13948e-39 = -8.74996e-39
	(b"00000000000100110100100100111011", b"00000000000000000000000000000000"),
	(b"00000000001011100010011010111011", b"00000000010000010110111111110110"), -- 1.77114e-39 + 4.23833e-39 = 6.00947e-39
	(b"00000000000011101101101101011101", b"00000000000000000000000000000000"),
	(b"00000000011000100011010100101000", b"00000000011100010001000010000101"), -- 1.36439e-39 + 9.01895e-39 = 1.03833e-38
	(b"10000000001001101110010001101001", b"00000000000000000000000000000000"),
	(b"00000000001011111111101010000110", b"00000000000010010001011000011101"), -- -3.57169e-39 + 4.40614e-39 = 8.34452e-40
	(b"00000000010011100101011001010010", b"00000000000000000000000000000000"),
	(b"10000000000011100111111101110111", b"00000000001111111101011011011011"), -- 7.19413e-39 + -1.33142e-39 = 5.86271e-39
	(b"10000000011000001000111000000101", b"00000000000000000000000000000000"),
	(b"00000000001001101000101110100011", b"10000000001110100000001001100010"), -- -8.86715e-39 + 3.53984e-39 = -5.32731e-39
	(b"00000000000001101101100100011110", b"00000000000000000000000000000000"),
	(b"00000000011111111111010111010010", b"00000000100001101100111011110000"), -- 6.289e-40 + 1.17513e-38 = 1.23802e-38
	(b"00000000010111110100010100001111", b"00000000000000000000000000000000"),
	(b"10000000010001110101111111001000", b"00000000000101111110010101000111"), -- 8.74915e-39 + -6.55468e-39 = 2.19447e-39
	(b"00000000001010101101100011110010", b"00000000000000000000000000000000"),
	(b"00000000011011110010101110011111", b"00000000100110100000010010010001"), -- 3.93492e-39 + 1.02094e-38 = 1.41443e-38
	(b"10000000011000101100100100001111", b"00000000000000000000000000000000"),
	(b"00000000011000110101111011000101", b"00000000000000001001010110110110"), -- -9.072e-39 + 9.12571e-39 = 5.37062e-41
	(b"10000000001101101010110100111001", b"00000000000000000000000000000000"),
	(b"10000000010011011100110011101000", b"10000000100001000111101000100001"), -- -5.02126e-39 + -7.14484e-39 = -1.21661e-38
	(b"10000000011011100000010001000110", b"00000000000000000000000000000000"),
	(b"10000000010110110110011100110000", b"10000000110010010110101101110110"), -- -1.01034e-38 + -8.39405e-39 = -1.84975e-38
	(b"00000000001001111100001000011010", b"00000000000000000000000000000000"),
	(b"10000000010101110101001011010000", b"10000000001011111001000010110110"), -- 3.65121e-39 + -8.0194e-39 = -4.36818e-39
	(b"00000000010001000101010010110111", b"00000000000000000000000000000000"),
	(b"00000000011111100001000111110011", b"00000000110000100110011010101010"), -- 6.2752e-39 + 1.15777e-38 = 1.78529e-38
	(b"00000000011001101100111010010111", b"00000000000000000000000000000000"),
	(b"00000000000111111010010101001001", b"00000000100001100111001111100000"), -- 9.44133e-39 + 2.90619e-39 = 1.23475e-38
	(b"00000000010111111110101011001110", b"00000000000000000000000000000000"),
	(b"10000000010110101101010110000000", b"00000000000001010001010101001110"), -- 8.8086e-39 + -8.34178e-39 = 4.6682e-40
	(b"10000000000101111000100111000000", b"00000000000000000000000000000000"),
	(b"10000000010000111011110100011010", b"10000000010110110100011011011010"), -- -2.16163e-39 + -6.22082e-39 = -8.38245e-39
	(b"00000000011010110110100010110000", b"00000000000000000000000000000000"),
	(b"00000000011010101001100011001110", b"00000000110101100000000101111110"), -- 9.86395e-39 + 9.78938e-39 = 1.96533e-38
	(b"10000000000110101011111001101100", b"00000000000000000000000000000000"),
	(b"10000000010011010000110111111110", b"10000000011001111100110001101010"), -- -2.45603e-39 + -7.07635e-39 = -9.53239e-39
	(b"10000000000110111110010110111000", b"00000000000000000000000000000000"),
	(b"00000000011101111111111110110010", b"00000000010111000001100111111010"), -- -2.56197e-39 + 1.10202e-38 = 8.45818e-39
	(b"10000000001101100101100001100001", b"00000000000000000000000000000000"),
	(b"10000000010111001010101101110110", b"10000000100100110000001111010111"), -- -4.99082e-39 + -8.51037e-39 = -1.35012e-38
	(b"10000000000011110100010100001000", b"00000000000000000000000000000000"),
	(b"00000000001111100101100001110010", b"00000000001011110001001101101010"), -- -1.4023e-39 + 5.72553e-39 = 4.32323e-39
	(b"00000000011111001111010100110111", b"00000000000000000000000000000000"),
	(b"10000000000110100101011111000101", b"00000000011000101001110101110010"), -- 1.14756e-38 + -2.41921e-39 = 9.05636e-39
	(b"10000000010100011101110001000110", b"00000000000000000000000000000000"),
	(b"10000000001011101100010101100010", b"10000000100000001010000110101000"), -- -7.51769e-39 + -4.29524e-39 = -1.18129e-38
	(b"10000000011101001111100100001010", b"00000000000000000000000000000000"),
	(b"10000000011000110000110000110100", b"10000000110110000000010100111110"), -- -1.07423e-38 + -9.09609e-39 = -1.98383e-38
	(b"00000000010010100101010111001100", b"00000000000000000000000000000000"),
	(b"10000000011010101110111001000101", b"10000000001000001001100001111001"), -- 6.8266e-39 + -9.82004e-39 = -2.99343e-39
	(b"00000000011010011111011111000100", b"00000000000000000000000000000000"),
	(b"00000000000010000000101001000000", b"00000000011100100000001000000100"), -- 9.73161e-39 + 7.38361e-40 = 1.047e-38
	(b"00000000011011101101000111100010", b"00000000000000000000000000000000"),
	(b"10000000001110111010101100100100", b"00000000001100110010011010111110"), -- 1.01772e-38 + -5.47969e-39 = 4.69751e-39
	(b"00000000000010111000101001101011", b"00000000000000000000000000000000"),
	(b"00000000000001101011010011111011", b"00000000000100100011111101100110"), -- 1.05985e-39 + 6.15937e-40 = 1.67578e-39
	(b"00000000011011110110100100001111", b"00000000000000000000000000000000"),
	(b"00000000010100100110000000101100", b"00000000110000011100100100111011"), -- 1.02314e-38 + 7.56501e-39 = 1.77964e-38
	(b"10000000001011001101101001110111", b"00000000000000000000000000000000"),
	(b"00000000001110011011000101110010", b"00000000000011001101011011111011"), -- -4.11913e-39 + 5.29828e-39 = 1.17915e-39
	(b"00000000001100011110010011000000", b"00000000000000000000000000000000"),
	(b"10000000010010111100100000000100", b"10000000000110011110001101000100"), -- 4.582e-39 + -6.95941e-39 = -2.37741e-39
	(b"10000000011001110110101110011100", b"00000000000000000000000000000000"),
	(b"00000000011111101110100010101000", b"00000000000101110111110100001100"), -- -9.49766e-39 + 1.16547e-38 = 2.15707e-39
	(b"10000000001000010000101101111001", b"00000000000000000000000000000000"),
	(b"00000000011001001111110101010101", b"00000000010000111111000111011100"), -- -3.03469e-39 + 9.27443e-39 = 6.23974e-39
	(b"00000000000101100111110100100100", b"00000000000000000000000000000000"),
	(b"10000000000000010101011010001011", b"00000000000101010010011010011001"), -- 2.06527e-39 + -1.22881e-40 = 1.94239e-39
	(b"00000000001101011001010111110101", b"00000000000000000000000000000000"),
	(b"00000000000100011000110010001101", b"00000000010001110010001010000010"), -- 4.92108e-39 + 1.61162e-39 = 6.5327e-39
	(b"10000000011001001101111100111101", b"00000000000000000000000000000000"),
	(b"00000000001100101010011101011010", b"10000000001100100011011111100011"), -- -9.26363e-39 + 4.65181e-39 = -4.61182e-39
	(b"10000000001001101001010001011100", b"00000000000000000000000000000000"),
	(b"00000000010001101111111100110100", b"00000000001000000110101011011000"), -- -3.54297e-39 + 6.52003e-39 = 2.97706e-39
	(b"10000000001001110101010000010011", b"00000000000000000000000000000000"),
	(b"10000000001000110111000001100001", b"10000000010010101100010001110100"), -- -3.61174e-39 + -3.25456e-39 = -6.8663e-39
	(b"00000000010100111011000011111111", b"00000000000000000000000000000000"),
	(b"00000000000110110010011011011100", b"00000000011011101101011111011011"), -- 7.68584e-39 + 2.4935e-39 = 1.01793e-38
	(b"00000000001000001110100010110011", b"00000000000000000000000000000000"),
	(b"10000000011100110000110010011100", b"10000000010100100010001111101001"), -- 3.02221e-39 + -1.05656e-38 = -7.54339e-39
	(b"00000000000110001010100100101100", b"00000000000000000000000000000000"),
	(b"10000000011100001010110000100001", b"10000000010110000000001011110101"), -- 2.26474e-39 + -1.03473e-38 = -8.08258e-39
	(b"10000000010010001011101001111010", b"00000000000000000000000000000000"),
	(b"10000000000010100000010101001101", b"10000000010100101011111111000111"), -- -6.67905e-39 + -9.20257e-40 = -7.59931e-39
	(b"10000000001100101100111000000011", b"00000000000000000000000000000000"),
	(b"10000000001000001101000110101011", b"10000000010100111001111110101110"), -- -4.66568e-39 + -3.01395e-39 = -7.67963e-39
	(b"00000000001001100001010010010011", b"00000000000000000000000000000000"),
	(b"10000000001100100000100111100011", b"10000000000010111111010101010000"), -- 3.49713e-39 + -4.59532e-39 = -1.09819e-39
	(b"00000000000111111100111000000111", b"00000000000000000000000000000000"),
	(b"00000000000101001011010100010011", b"00000000001101001000001100011010"), -- 2.92081e-39 + 1.90167e-39 = 4.82248e-39
	(b"10000000011101100110100100001110", b"00000000000000000000000000000000"),
	(b"00000000001101110001110101010000", b"10000000001111110100101110111110"), -- -1.08743e-38 + 5.06147e-39 = -5.81281e-39
	(b"10000000001000000101111111001110", b"00000000000000000000000000000000"),
	(b"10000000001001111101001011100101", b"10000000010010000011001010110011"), -- -2.9731e-39 + -3.65724e-39 = -6.63034e-39
	(b"10000000001010011010011000111111", b"00000000000000000000000000000000"),
	(b"00000000010011100000001010001110", b"00000000001001000101110001001111"), -- -3.82489e-39 + 7.16409e-39 = 3.33919e-39
	(b"10000000011111110101100011000100", b"00000000000000000000000000000000"),
	(b"00000000010011110001011010010001", b"10000000001100000100001000110011"), -- -1.1695e-38 + 7.2631e-39 = -4.43185e-39
	(b"00000000001101101010010011011111", b"00000000000000000000000000000000"),
	(b"00000000011110011100000000001111", b"00000000101100000110010011101110"), -- 5.01826e-39 + 1.1181e-38 = 1.61993e-38
	(b"10000000001011110001001110110110", b"00000000000000000000000000000000"),
	(b"10000000001001010101101011101111", b"10000000010101000110111010100101"), -- -4.32334e-39 + -3.43053e-39 = -7.75387e-39
	(b"00000000010011011010111110001101", b"00000000000000000000000000000000"),
	(b"00000000011100001100000100101001", b"00000000101111100111000010110110"), -- 7.13431e-39 + 1.03549e-38 = 1.74892e-38
	(b"10000000010001001010010001110011", b"00000000000000000000000000000000"),
	(b"00000000011111110111100001000111", b"00000000001110101101001111010100"), -- -6.30381e-39 + 1.17063e-38 = 5.40245e-39
	(b"00000000011000111110111001111001", b"00000000000000000000000000000000"),
	(b"00000000001011011101100100101000", b"00000000100100011100011110100001"), -- 9.17726e-39 + 4.2105e-39 = 1.33878e-38
	(b"00000000010001110110111010000111", b"00000000000000000000000000000000"),
	(b"10000000010011001001000001010000", b"10000000000001010010000111001001"), -- 6.55997e-39 + -7.03127e-39 = -4.71297e-40
	(b"00000000001001000101100110100100", b"00000000000000000000000000000000"),
	(b"10000000010001001101111000100000", b"10000000001000001000010001111100"), -- 3.33823e-39 + -6.3245e-39 = -2.98626e-39
	(b"10000000010010101011100110000000", b"00000000000000000000000000000000"),
	(b"00000000011011110111111000011101", b"00000000001001001100010010011101"), -- -6.86237e-39 + 1.0239e-38 = 3.37661e-39
	(b"10000000010000100100100000101001", b"00000000000000000000000000000000"),
	(b"00000000011110010011010110011011", b"00000000001101101110110101110010"), -- -6.08703e-39 + 1.11313e-38 = 5.0443e-39
	(b"10000000010100100000110000001110", b"00000000000000000000000000000000"),
	(b"10000000000110101011011011110001", b"10000000011011001100001011111111"), -- -7.53484e-39 + -2.45335e-39 = -9.98819e-39
	(b"00000000010100000010000000101111", b"00000000000000000000000000000000"),
	(b"00000000000001001100010011010010", b"00000000010101001110010100000001"), -- 7.35838e-39 + 4.37948e-40 = 7.79633e-39
	(b"10000000000110010000111100001100", b"00000000000000000000000000000000"),
	(b"10000000000101111110101001100100", b"10000000001100001111100101110000"), -- -2.30129e-39 + -2.1963e-39 = -4.49759e-39
	(b"10000000011110011011001001001100", b"00000000000000000000000000000000"),
	(b"10000000010101001001000001111000", b"10000000110011100100001011000100"), -- -1.11761e-38 + -7.76601e-39 = -1.89421e-38
	(b"00000000011110111101001110001010", b"00000000000000000000000000000000"),
	(b"10000000011010101101001100010001", b"00000000000100010000000001111001"), -- 1.13717e-38 + -9.81028e-39 = 1.56137e-39
	(b"00000000001101100010101001010111", b"00000000000000000000000000000000"),
	(b"00000000010100101010001110101110", b"00000000100010001100111000000101"), -- 4.97431e-39 + 7.58923e-39 = 1.25635e-38
	(b"00000000000000010001001100011100", b"00000000000000000000000000000000"),
	(b"00000000000111011100001111111110", b"00000000000111101101011100011010"), -- 9.86906e-41 + 2.73354e-39 = 2.83223e-39
	(b"10000000000000011010010101110111", b"00000000000000000000000000000000"),
	(b"00000000011110000010101110110101", b"00000000011101101000011000111110"), -- -1.51193e-40 + 1.10359e-38 = 1.08847e-38
	(b"10000000001100110011100011001011", b"00000000000000000000000000000000"),
	(b"10000000001011010111000100100111", b"10000000011000001010100111110010"), -- -4.70398e-39 + -4.17319e-39 = -8.87717e-39
	(b"00000000011000110000010111010100", b"00000000000000000000000000000000"),
	(b"10000000011101001101100011100100", b"10000000000100011101001100010000"), -- 9.0938e-39 + -1.07307e-38 = -1.63692e-39
	(b"10000000010001100011000100011000", b"00000000000000000000000000000000"),
	(b"00000000000111101011111100010111", b"10000000001001110111001000000001"), -- -6.4461e-39 + 2.82362e-39 = -3.62248e-39
	(b"10000000010100101111000000000011", b"00000000000000000000000000000000"),
	(b"00000000001010011110111110000111", b"10000000001010010000000001111100"), -- -7.61661e-39 + 3.85118e-39 = -3.76543e-39
	(b"00000000011110101110110011011000", b"00000000000000000000000000000000"),
	(b"10000000001101100100011100010001", b"00000000010001001010010111000111"), -- 1.12889e-38 + -4.98461e-39 = 6.30428e-39
	(b"10000000000110001110010000110111", b"00000000000000000000000000000000"),
	(b"00000000001010001010100100101101", b"00000000000011111100010011110110"), -- -2.28592e-39 + 3.73411e-39 = 1.44819e-39
	(b"00000000001111100110010011011000", b"00000000000000000000000000000000"),
	(b"00000000010010011100001001110110", b"00000000100010000010011101001110"), -- 5.72998e-39 + 6.77375e-39 = 1.25037e-38
	(b"00000000011011100100100101110110", b"00000000000000000000000000000000"),
	(b"00000000010101101000000100110110", b"00000000110001001100101010101100"), -- 1.01283e-38 + 7.9442e-39 = 1.80725e-38
	(b"10000000000000000100111000100001", b"00000000000000000000000000000000"),
	(b"10000000000110111111000100000010", b"10000000000111000011111100100011"), -- -2.80274e-41 + -2.56602e-39 = -2.59404e-39
	(b"00000000010101011110110010110100", b"00000000000000000000000000000000"),
	(b"00000000001111111111010110100101", b"00000000100101011110001001011001"), -- 7.89093e-39 + 5.87376e-39 = 1.37647e-38
	(b"00000000010001101110000101011010", b"00000000000000000000000000000000"),
	(b"00000000001010011010111100101011", b"00000000011100001001000010000101"), -- 6.50933e-39 + 3.82809e-39 = 1.03374e-38
	(b"10000000000011010100000010001000", b"00000000000000000000000000000000"),
	(b"00000000001111100100000011011011", b"00000000001100010000000001010011"), -- -1.21701e-39 + 5.71707e-39 = 4.50006e-39
	(b"10000000000000001100101110000010", b"00000000000000000000000000000000"),
	(b"00000000011101101001111011010001", b"00000000011101011101001101001111"), -- -7.30048e-41 + 1.08936e-38 = 1.08206e-38
	(b"00000000001100010100110111110101", b"00000000000000000000000000000000"),
	(b"00000000000011100001110101100011", b"00000000001111110110101101011000"), -- 4.52791e-39 + 1.29624e-39 = 5.82414e-39
	(b"10000000010011101001011010010010", b"00000000000000000000000000000000"),
	(b"10000000010110001001001010000100", b"10000000101001110010100100010110"), -- -7.21718e-39 + -8.13408e-39 = -1.53513e-38
	(b"00000000010010001110010100010111", b"00000000000000000000000000000000"),
	(b"00000000000011000001000110000111", b"00000000010101001111011010011110"), -- 6.69434e-39 + 1.10831e-39 = 7.80265e-39
	(b"00000000000110111010001101100011", b"00000000000000000000000000000000"),
	(b"00000000000011101000101110001111", b"00000000001010100010111011110010"), -- 2.53817e-39 + 1.33576e-39 = 3.87393e-39
	(b"10000000011111000000000111010110", b"00000000000000000000000000000000"),
	(b"10000000001010001110100010001110", b"10000000101001001110101001100100"), -- -1.13883e-38 + -3.75684e-39 = -1.51451e-38
	(b"10000000011101100110001111101110", b"00000000000000000000000000000000"),
	(b"00000000001100011000010101011010", b"10000000010001001101111010010100"), -- -1.08724e-38 + 4.54778e-39 = -6.32466e-39
	(b"10000000000000011101101000011111", b"00000000000000000000000000000000"),
	(b"10000000010101010001000111011010", b"10000000010101101110101111111001"), -- -1.70083e-40 + -7.81242e-39 = -7.9825e-39
	(b"10000000000010101000110010011010", b"00000000000000000000000000000000"),
	(b"00000000010111100000110110001101", b"00000000010100111000000011110011"), -- -9.68793e-40 + 8.6374e-39 = 7.6686e-39
	(b"00000000000011100111001010111010", b"00000000000000000000000000000000"),
	(b"00000000000110100011011001011000", b"00000000001010001010100100010010"), -- 1.32685e-39 + 2.40722e-39 = 3.73407e-39
	(b"10000000001001010001001101001001", b"00000000000000000000000000000000"),
	(b"10000000001011101101110101110110", b"10000000010100111111000010111111"), -- -3.40483e-39 + -4.30388e-39 = -7.70871e-39
	(b"10000000000100001110100111000001", b"00000000000000000000000000000000"),
	(b"00000000000101011000011100110001", b"00000000000001001001110101110000"), -- -1.55322e-39 + 1.97704e-39 = 4.2382e-40
	(b"00000000000010110001101111011011", b"00000000000000000000000000000000"),
	(b"00000000000000101101001001100010", b"00000000000011011110111000111101"), -- 1.02018e-39 + 2.59142e-40 = 1.27933e-39
	(b"10000000010011100001101000010001", b"00000000000000000000000000000000"),
	(b"10000000001010001010111101111010", b"10000000011101101100100110001011"), -- -7.17252e-39 + -3.73637e-39 = -1.09089e-38
	(b"00000000000111100001110101000000", b"00000000000000000000000000000000"),
	(b"00000000000110111101011110000010", b"00000000001110011111010011000010"), -- 2.76556e-39 + 2.55687e-39 = 5.32243e-39
	(b"00000000000111100011001001010010", b"00000000000000000000000000000000"),
	(b"10000000010001101001000111110110", b"10000000001010000101111110100100"), -- 2.77312e-39 + -6.48085e-39 = -3.70773e-39
	(b"10000000001010001011011100101011", b"00000000000000000000000000000000"),
	(b"00000000010001110011000111010010", b"00000000000111100111101010100111"), -- -3.73913e-39 + 6.53819e-39 = 2.79906e-39
	(b"10000000010001001110000010010011", b"00000000000000000000000000000000"),
	(b"10000000011101110100110110100011", b"10000000101111000010111000110110"), -- -6.32538e-39 + -1.09563e-38 = -1.72817e-38
	(b"10000000011110011111010010110101", b"00000000000000000000000000000000"),
	(b"00000000000010101000110101111010", b"10000000011011110110011100111011"), -- -1.11999e-38 + 9.69107e-40 = -1.02308e-38
	(b"00000000010011101110101101111010", b"00000000000000000000000000000000"),
	(b"00000000001100001100001001010010", b"00000000011111111010110111001100"), -- 7.24764e-39 + 4.47781e-39 = 1.17255e-38
	(b"00000000010100101010001110011001", b"00000000000000000000000000000000"),
	(b"10000000001110000011010010010000", b"00000000000110100110111100001001"), -- 7.5892e-39 + -5.16164e-39 = 2.42755e-39
	(b"00000000011011001011101111101001", b"00000000000000000000000000000000"),
	(b"10000000000111011111100000011110", b"00000000010011101100001111001011"), -- 9.98564e-39 + -2.75224e-39 = 7.23341e-39
	(b"10000000010110101110000111111110", b"00000000000000000000000000000000"),
	(b"00000000001110000000011100011100", b"10000000001000101101101011100010"), -- -8.34627e-39 + 5.14534e-39 = -3.20093e-39
	(b"10000000010101111110000101011101", b"00000000000000000000000000000000"),
	(b"10000000010101110001100000111110", b"10000000101011101111100110011011"), -- -8.07053e-39 + -7.99838e-39 = -1.60689e-38
	(b"10000000010110111011101100011011", b"00000000000000000000000000000000"),
	(b"00000000011111111010000111011001", b"00000000001000111110011010111110"), -- -8.42415e-39 + 1.17212e-38 = 3.29702e-39
	(b"10000000001101110111100110011010", b"00000000000000000000000000000000"),
	(b"10000000010101110110111001010011", b"10000000100011101110011111101101"), -- -5.09457e-39 + -8.02927e-39 = -1.31238e-38
	(b"00000000000000100111100100100010", b"00000000000000000000000000000000"),
	(b"10000000011110010111000110011011", b"10000000011101101111100001111001"), -- 2.27125e-40 + -1.11528e-38 = -1.09257e-38
	(b"00000000010000010111011001101000", b"00000000000000000000000000000000"),
	(b"10000000000000001100111110000001", b"00000000010000001010011011100111"), -- 6.01178e-39 + -7.44384e-41 = 5.93735e-39
	(b"10000000010110011111010001011001", b"00000000000000000000000000000000"),
	(b"10000000001011100110111110010000", b"10000000100010000110001111101001"), -- -8.26101e-39 + -4.26445e-39 = -1.25255e-38
	(b"00000000001100010111010001011010", b"00000000000000000000000000000000"),
	(b"00000000010101100100000011001011", b"00000000100001111011010100100101"), -- 4.54168e-39 + 7.9211e-39 = 1.24628e-38
	(b"10000000010001111111100111010001", b"00000000000000000000000000000000"),
	(b"00000000010100001111101101001111", b"00000000000010010000000101111110"), -- -6.60994e-39 + 7.43699e-39 = 8.27055e-40
	(b"10000000010000010011001011000110", b"00000000000000000000000000000000"),
	(b"00000000000011011101000111000000", b"10000000001100110110000100000110"), -- -5.98752e-39 + 1.26911e-39 = -4.71842e-39
	(b"10000000000110101001010110010110", b"00000000000000000000000000000000"),
	(b"00000000001100100100000001110100", b"00000000000101111010101011011110"), -- -2.44138e-39 + 4.6149e-39 = 2.17351e-39
	(b"10000000010111011110101010111100", b"00000000000000000000000000000000"),
	(b"00000000000011010100000010111100", b"10000000010100001010101000000000"), -- -8.62491e-39 + 1.21708e-39 = -7.40782e-39
	(b"00000000010100100111110011100010", b"00000000000000000000000000000000"),
	(b"10000000010010011110010010011110", b"00000000000010001001100001000100"), -- 7.57531e-39 + -6.786e-39 = 7.89307e-40
	(b"10000000011001111001111001100110", b"00000000000000000000000000000000"),
	(b"10000000010010100111001011001101", b"10000000101100100001000100110011"), -- -9.51588e-39 + -6.83701e-39 = -1.63529e-38
	(b"10000000010001100111001111011110", b"00000000000000000000000000000000"),
	(b"10000000000110000010101100011110", b"10000000010111101001111011111100"), -- -6.47005e-39 + -2.21952e-39 = -8.68957e-39
	(b"10000000001101101100110110010111", b"00000000000000000000000000000000"),
	(b"00000000001111000010000100001001", b"00000000000001010101001101110010"), -- -5.03287e-39 + 5.52198e-39 = 4.89112e-40
	(b"00000000001101001011010101101010", b"00000000000000000000000000000000"),
	(b"10000000001001001111100011001011", b"00000000000011111011110010011111"), -- 4.84052e-39 + -3.39533e-39 = 1.4452e-39
	(b"00000000011100100001000010000000", b"00000000000000000000000000000000"),
	(b"00000000000001011100010000101000", b"00000000011101111101010010101000"), -- 1.04752e-38 + 5.29545e-40 = 1.10047e-38
	(b"00000000011101110011001111001010", b"00000000000000000000000000000000"),
	(b"00000000000001111001110011110010", b"00000000011111101101000010111100"), -- 1.0947e-38 + 6.9915e-40 = 1.16462e-38
	(b"00000000000110101000100110010010", b"00000000000000000000000000000000"),
	(b"00000000001011101010010011111011", b"00000000010010010010111010001101"), -- 2.43707e-39 + 4.28362e-39 = 6.72069e-39
	(b"00000000010100001110011100011101", b"00000000000000000000000000000000"),
	(b"00000000011110000100100010110111", b"00000000110010010010111111010100"), -- 7.42975e-39 + 1.10463e-38 = 1.84761e-38
	(b"10000000010001101000011001000111", b"00000000000000000000000000000000"),
	(b"00000000000111110010110101101101", b"10000000001001110101100011011010"), -- -6.47665e-39 + 2.8632e-39 = -3.61346e-39
	(b"10000000001110001001010100011010", b"00000000000000000000000000000000"),
	(b"10000000001110001110100010100000", b"10000000011100010111110110111010"), -- -5.19628e-39 + -5.22624e-39 = -1.04225e-38
	(b"10000000011011100000011101001001", b"00000000000000000000000000000000"),
	(b"00000000000001010111000110011101", b"10000000011010001001010110101100"), -- -1.01045e-38 + 4.99934e-40 = -9.60458e-39
	(b"00000000001001100111110111100111", b"00000000000000000000000000000000"),
	(b"00000000001110101010110111010011", b"00000000011000010010101110111010"), -- 3.53491e-39 + 5.38882e-39 = 8.92373e-39
	(b"00000000010101100000110111110000", b"00000000000000000000000000000000"),
	(b"00000000001100000001110010100110", b"00000000100001100010101010010110"), -- 7.90285e-39 + 4.41838e-39 = 1.23212e-38
	(b"10000000011001010000000100011000", b"00000000000000000000000000000000"),
	(b"00000000000000111011000100111100", b"10000000011000010100111111011100"), -- -9.27578e-39 + 3.39086e-40 = -8.93669e-39
	(b"10000000001001000101100000101110", b"00000000000000000000000000000000"),
	(b"00000000010011110110010010111000", b"00000000001010110000110010001010"), -- -3.33771e-39 + 7.29114e-39 = 3.95342e-39
	(b"00000000000101111000001000111010", b"00000000000000000000000000000000"),
	(b"00000000010110110111011010010001", b"00000000011100101111100011001011"), -- 2.15893e-39 + 8.39956e-39 = 1.05585e-38
	(b"00000000010011111100010100100100", b"00000000000000000000000000000000"),
	(b"10000000000110101010110110111010", b"00000000001101010001011101101010"), -- 7.32572e-39 + -2.45004e-39 = 4.87568e-39
	(b"00000000000010111000000111010101", b"00000000000000000000000000000000"),
	(b"00000000000101011010111110110000", b"00000000001000010011000110000101"), -- 1.05677e-39 + 1.99157e-39 = 3.04834e-39
	(b"10000000010100101110101000101010", b"00000000000000000000000000000000"),
	(b"10000000010001110100010011000011", b"10000000100110100010111011101101"), -- -7.61451e-39 + -6.54499e-39 = -1.41595e-38
	(b"10000000011110110101011111011000", b"00000000000000000000000000000000"),
	(b"10000000001111110100011000101110", b"10000000101110101001111000000110"), -- -1.13273e-38 + -5.81081e-39 = -1.71381e-38
	(b"00000000000010101101100101111011", b"00000000000000000000000000000000"),
	(b"10000000010101010000000001101000", b"10000000010010100010011011101101"), -- 9.96372e-40 + -7.80616e-39 = -6.80979e-39
	(b"00000000011010000000101100000011", b"00000000000000000000000000000000"),
	(b"00000000001100010111110000001111", b"00000000100110011000011100010010"), -- 9.55484e-39 + 4.54444e-39 = 1.40993e-38
	(b"00000000011001011000000011000100", b"00000000000000000000000000000000"),
	(b"10000000010011010111100101101111", b"00000000000110000000011101010101"), -- 9.32158e-39 + -7.1149e-39 = 2.20668e-39
	(b"10000000011001000100110100101000", b"00000000000000000000000000000000"),
	(b"10000000011110011010001000001101", b"10000000110111011110111100110101"), -- -9.21123e-39 + -1.11702e-38 = -2.03815e-38
	(b"00000000001101001010101001000011", b"00000000000000000000000000000000"),
	(b"00000000001010000010001100111011", b"00000000010111001100110101111110"), -- 4.83652e-39 + 3.68606e-39 = 8.52258e-39
	(b"10000000010011111010101110011100", b"00000000000000000000000000000000"),
	(b"00000000001110101100001011001000", b"10000000000101001110100011010100"), -- -7.31657e-39 + 5.39633e-39 = -1.92023e-39
	(b"10000000000111000000100011000110", b"00000000000000000000000000000000"),
	(b"00000000010110100010000111000011", b"00000000001111100001100011111101"), -- -2.57454e-39 + 8.27731e-39 = 5.70276e-39
	(b"10000000001010010111100100100111", b"00000000000000000000000000000000"),
	(b"10000000001110100011101110100110", b"10000000011000111011010011001101"), -- -3.80872e-39 + -5.34786e-39 = -9.15657e-39
	(b"00000000010000000111100111010010", b"00000000000000000000000000000000"),
	(b"10000000000001111001011111101100", b"00000000001110001110000111100110"), -- 5.92117e-39 + -6.97348e-40 = 5.22382e-39
	(b"00000000011101001001111001100010", b"00000000000000000000000000000000"),
	(b"10000000001000110011000110001101", b"00000000010100010110110011010101"), -- 1.07097e-38 + -3.23202e-39 = 7.47772e-39
	(b"00000000000110100011001110001111", b"00000000000000000000000000000000"),
	(b"10000000010001010010111011001100", b"10000000001010101111101100111101"), -- 2.40622e-39 + -6.35344e-39 = -3.94722e-39
	(b"00000000000000111001010110110001", b"00000000000000000000000000000000"),
	(b"00000000000101111001000101100010", b"00000000000110110010011100010011"), -- 3.29206e-40 + 2.16437e-39 = 2.49358e-39
	(b"00000000001001111110101101111110", b"00000000000000000000000000000000"),
	(b"00000000000101111101000111100000", b"00000000001111111011110101011110"), -- 3.66606e-39 + 2.18751e-39 = 5.85357e-39
	(b"00000000001011111101010110101011", b"00000000000000000000000000000000"),
	(b"00000000000100010100001101001011", b"00000000010000010001100011110110"), -- 4.39292e-39 + 1.58534e-39 = 5.97826e-39
	(b"00000000010010001100111010011011", b"00000000000000000000000000000000"),
	(b"00000000010101101111011011110000", b"00000000100111111100010110001011"), -- 6.68627e-39 + 7.98644e-39 = 1.46727e-38
	(b"10000000010110000110111100110000", b"00000000000000000000000000000000"),
	(b"10000000011010101110101101010101", b"10000000110000110101101010000101"), -- -8.12141e-39 + -9.81898e-39 = -1.79404e-38
	(b"10000000010011101000100001010001", b"00000000000000000000000000000000"),
	(b"00000000001110110000101011110110", b"10000000000100110111110101011011"), -- -7.21207e-39 + 5.42223e-39 = -1.78984e-39
	(b"00000000010011010000101011010001", b"00000000000000000000000000000000"),
	(b"10000000000000001000100000010000", b"00000000010011001000001011000001"), -- 7.07521e-39 + -4.881e-41 = 7.0264e-39
	(b"00000000001101000000111101011010", b"00000000000000000000000000000000"),
	(b"00000000010010101001100011110111", b"00000000011111101010100001010001"), -- 4.78095e-39 + 6.8507e-39 = 1.16317e-38
	(b"10000000010111000111111000100011", b"00000000000000000000000000000000"),
	(b"00000000001011011010110000000100", b"10000000001011101101001000011111"), -- -8.49411e-39 + 4.1943e-39 = -4.29981e-39
	(b"10000000011000111011101111011011", b"00000000000000000000000000000000"),
	(b"10000000010011010111011101111001", b"10000000101100010011001101010100"), -- -9.1591e-39 + -7.11419e-39 = -1.62733e-38
	(b"00000000001011011110100110110111", b"00000000000000000000000000000000"),
	(b"00000000001011000010001000111000", b"00000000010110100000101111101111"), -- 4.21644e-39 + 4.05304e-39 = 8.26948e-39
	(b"00000000011110001100100101011001", b"00000000000000000000000000000000"),
	(b"00000000010101111110011111010101", b"00000000110100001011000100101110"), -- 1.10925e-38 + 8.07285e-39 = 1.91653e-38
	(b"00000000001001110000010010100110", b"00000000000000000000000000000000"),
	(b"10000000010101010010000000000111", b"10000000001011100001101101100001"), -- 3.58325e-39 + -7.81751e-39 = -4.23425e-39
	(b"00000000010010001111110110001000", b"00000000000000000000000000000000"),
	(b"00000000010000110011100000000011", b"00000000100011000011010110001011"), -- 6.70311e-39 + 6.17307e-39 = 1.28762e-38
	(b"10000000010010010001110111111010", b"00000000000000000000000000000000"),
	(b"10000000001110101011110100111011", b"10000000100000111101101100110101"), -- -6.71474e-39 + -5.39434e-39 = -1.21091e-38
	(b"10000000001001011010010111000010", b"00000000000000000000000000000000"),
	(b"00000000010110111011011010110101", b"00000000001101100001000011110011"), -- -3.45738e-39 + 8.42257e-39 = 4.9652e-39
	(b"10000000011111101111101001000100", b"00000000000000000000000000000000"),
	(b"10000000001011010011010011100100", b"10000000101011000010111100101000"), -- -1.16611e-38 + -4.15157e-39 = -1.58126e-38
	(b"00000000000111000011000001110010", b"00000000000000000000000000000000"),
	(b"10000000010001111100010010000111", b"10000000001010111001010000010101"), -- 2.58877e-39 + -6.59082e-39 = -4.00205e-39
	(b"00000000001100001100010111111001", b"00000000000000000000000000000000"),
	(b"00000000011111111010001010000001", b"00000000101100000110100001111010"), -- 4.47912e-39 + 1.17214e-38 = 1.62005e-38
	(b"10000000010100000010001101100001", b"00000000000000000000000000000000"),
	(b"10000000001011100010000111000001", b"10000000011111100100010100100010"), -- -7.35953e-39 + -4.23654e-39 = -1.15961e-38
	(b"10000000001110000000111100111100", b"00000000000000000000000000000000"),
	(b"00000000001010111100111111000111", b"10000000000011000011111101110101"), -- -5.14825e-39 + 4.02346e-39 = -1.12479e-39
	(b"10000000000001101010011001111111", b"00000000000000000000000000000000"),
	(b"00000000001110111110010101110000", b"00000000001101010011111011110001"), -- -6.10741e-40 + 5.5006e-39 = 4.88986e-39
	(b"00000000001110110010101001001011", b"00000000000000000000000000000000"),
	(b"00000000011111100010010110001000", b"00000000101110010100111111010011"), -- 5.43347e-39 + 1.15847e-38 = 1.70182e-38
	(b"10000000001000101000110101101001", b"00000000000000000000000000000000"),
	(b"10000000001001011011010100010010", b"10000000010010000100001001111011"), -- -3.17314e-39 + -3.46287e-39 = -6.636e-39
	(b"00000000000110011001110010111001", b"00000000000000000000000000000000"),
	(b"00000000010110001000010001101101", b"00000000011100100010000100100110"), -- 2.35211e-39 + 8.12903e-39 = 1.04811e-38
	(b"00000000010001000110001110000011", b"00000000000000000000000000000000"),
	(b"10000000000110001001111110010000", b"00000000001010111100001111110011"), -- 6.28051e-39 + -2.26129e-39 = 4.01922e-39
	(b"00000000010001000100111111000010", b"00000000000000000000000000000000"),
	(b"10000000011001111110011010100000", b"10000000001000111001011011011110"), -- 6.27343e-39 + -9.54179e-39 = -3.26836e-39
	(b"00000000010010100010010001001110", b"00000000000000000000000000000000"),
	(b"10000000000011101101100001110101", b"00000000001110110100101111011001"), -- 6.80885e-39 + -1.36335e-39 = 5.4455e-39
	(b"00000000000110111100001111111100", b"00000000000000000000000000000000"),
	(b"10000000011011011100100101001110", b"10000000010100100000010101010010"), -- 2.54986e-39 + -1.00823e-38 = -7.53242e-39
	(b"00000000001010111010101111001111", b"00000000000000000000000000000000"),
	(b"00000000001101110111001101111000", b"00000000011000110001111101000111"), -- 4.01056e-39 + 5.09237e-39 = 9.10293e-39
	(b"00000000001110000001011001001101", b"00000000000000000000000000000000"),
	(b"00000000000010010010110011100001", b"00000000010000010100001100101110"), -- 5.15079e-39 + 8.42619e-40 = 5.99341e-39
	(b"00000000010111011111000100000111", b"00000000000000000000000000000000"),
	(b"10000000010111010100000011100100", b"00000000000000001011000000100011"), -- 8.62717e-39 + -8.56398e-39 = 6.31859e-41
	(b"10000000001111100011001111000001", b"00000000000000000000000000000000"),
	(b"10000000000011101101101111001000", b"10000000010011010000111110001001"), -- -5.71237e-39 + -1.36454e-39 = -7.07691e-39
	(b"00000000000011110011000110101001", b"00000000000000000000000000000000"),
	(b"10000000010101000001111010001111", b"10000000010001001110110011100110"), -- 1.39535e-39 + -7.72514e-39 = -6.3298e-39
	(b"00000000010010110001101101110001", b"00000000000000000000000000000000"),
	(b"10000000001001111000110100000110", b"00000000001000111000111001101011"), -- 6.89751e-39 + -3.63217e-39 = 3.26533e-39
	(b"00000000010001101001110110000000", b"00000000000000000000000000000000"),
	(b"00000000011101001100101011100010", b"00000000101110110110100001100010"), -- 6.48499e-39 + 1.07257e-38 = 1.72107e-38
	(b"00000000010100101101011001000111", b"00000000000000000000000000000000"),
	(b"00000000000110101110010100101010", b"00000000011011011011101101110001"), -- 7.60738e-39 + 2.46993e-39 = 1.00773e-38
	(b"00000000001100011111110011100100", b"00000000000000000000000000000000"),
	(b"10000000011011110101001000001110", b"10000000001111010101010100101010"), -- 4.59066e-39 + -1.02232e-38 = -5.63252e-39
	(b"10000000010001111011000111101101", b"00000000000000000000000000000000"),
	(b"00000000001110100010100100011001", b"10000000000011011000100011010100"), -- -6.58415e-39 + 5.3412e-39 = -1.24295e-39
	(b"00000000010011100111110101000011", b"00000000000000000000000000000000"),
	(b"10000000000011111001100111101100", b"00000000001111101110001101010111"), -- 7.2081e-39 + -1.43275e-39 = 5.77535e-39
	(b"00000000011111111000001010010001", b"00000000000000000000000000000000"),
	(b"00000000001011101001001110101010", b"00000000101011100001011000111011"), -- 1.17099e-38 + 4.2774e-39 = 1.59874e-38
	(b"10000000011001110101100001101000", b"00000000000000000000000000000000"),
	(b"00000000001011010110010101100111", b"10000000001110011111001100000001"), -- -9.49077e-39 + 4.16897e-39 = -5.3218e-39
	(b"10000000010101001010101101001111", b"00000000000000000000000000000000"),
	(b"00000000001101101110101100110111", b"10000000000111011100000000011000"), -- -7.77564e-39 + 5.0435e-39 = -2.73214e-39
	(b"10000000010101011110100000100101", b"00000000000000000000000000000000"),
	(b"10000000001001111001010101101001", b"10000000011111010111110110001110"), -- -7.88929e-39 + -3.63518e-39 = -1.15245e-38
	(b"10000000000101010001111010101001", b"00000000000000000000000000000000"),
	(b"00000000000010111010010111100100", b"10000000000010010111100011000101"), -- -1.93954e-39 + 1.0697e-39 = -8.69843e-40
	(b"00000000000011111101101100010110", b"00000000000000000000000000000000"),
	(b"10000000010101010000001110000001", b"10000000010001010010100001101011"), -- 1.45613e-39 + -7.80727e-39 = -6.35115e-39
	(b"10000000001100011100100001110101", b"00000000000000000000000000000000"),
	(b"10000000010001110011110111101100", b"10000000011110010000011001100001"), -- -4.57185e-39 + -6.54253e-39 = -1.11144e-38
	(b"00000000000100111000001011000110", b"00000000000000000000000000000000"),
	(b"00000000000001111010110111011110", b"00000000000110110011000010100100"), -- 1.79179e-39 + 7.0522e-40 = 2.49701e-39
	(b"00000000001001111111001111000011", b"00000000000000000000000000000000"),
	(b"00000000001011000101010000011110", b"00000000010101000100011111100001"), -- 3.66903e-39 + 4.07094e-39 = 7.73997e-39
	(b"00000000000101100001000101011110", b"00000000000000000000000000000000"),
	(b"10000000011011011100011011000111", b"10000000010101111011010101101001"), -- 2.02661e-39 + -1.00814e-38 = -8.05477e-39
	(b"00000000000111110001010110001110", b"00000000000000000000000000000000"),
	(b"10000000011100100101110011010110", b"10000000010100110100011101001000"), -- 2.85463e-39 + -1.05025e-38 = -7.64792e-39
	(b"10000000001100010011100111110010", b"00000000000000000000000000000000"),
	(b"00000000001000001000110101101010", b"10000000000100001010110010001000"), -- -4.52073e-39 + 2.98947e-39 = -1.53126e-39
	(b"10000000011000111111100111010010", b"00000000000000000000000000000000"),
	(b"00000000001101001001100001010010", b"10000000001011110110000110000000"), -- -9.18133e-39 + 4.83009e-39 = -4.35124e-39
	(b"00000000011010110011101100110110", b"00000000000000000000000000000000"),
	(b"10000000000100011100010000101000", b"00000000010110010111011100001110"), -- 9.84764e-39 + -1.63157e-39 = 8.21607e-39
	(b"10000000001000010010011001000110", b"00000000000000000000000000000000"),
	(b"00000000011010101001101110010101", b"00000000010010010111010101001111"), -- -3.0443e-39 + 9.79037e-39 = 6.74607e-39
	(b"10000000010101011001011000001110", b"00000000000000000000000000000000"),
	(b"10000000011111011101110000110010", b"10000000110100110111001001000000"), -- -7.85985e-39 + -1.15584e-38 = -1.94183e-38
	(b"00000000001110111100110000101101", b"00000000000000000000000000000000"),
	(b"00000000011111111100100101111111", b"00000000101110111001010110101100"), -- 5.49154e-39 + 1.17354e-38 = 1.72269e-38
	(b"10000000001000111111110000001001", b"00000000000000000000000000000000"),
	(b"10000000010100110111011011110111", b"10000000011101110111001100000000"), -- -3.30466e-39 + -7.66502e-39 = -1.09697e-38
	(b"00000000010101010111011010010111", b"00000000000000000000000000000000"),
	(b"00000000001101100011000010001010", b"00000000100010111010011100100001"), -- 7.84856e-39 + 4.97653e-39 = 1.28251e-38
	(b"10000000000110110010101111101100", b"00000000000000000000000000000000"),
	(b"00000000001100001010110111011100", b"00000000000101011000000111110000"), -- -2.49531e-39 + 4.47047e-39 = 1.97516e-39
	(b"00000000011111011110101000111010", b"00000000000000000000000000000000"),
	(b"10000000001001001110111000011000", b"00000000010110001111110000100010"), -- 1.15635e-38 + -3.39149e-39 = 8.17197e-39
	(b"10000000001101111100101010100100", b"00000000000000000000000000000000"),
	(b"00000000011001010101110101100100", b"00000000001011011001001011000000"), -- -5.12365e-39 + 9.30889e-39 = 4.18524e-39
	(b"10000000000100010110110001001110", b"00000000000000000000000000000000"),
	(b"10000000010000110110100111000001", b"10000000010101001101011000001111"), -- -1.60006e-39 + -6.19092e-39 = -7.79097e-39
	(b"00000000010101110111100011101000", b"00000000000000000000000000000000"),
	(b"10000000011111111110101010100101", b"10000000001010000111000110111101"), -- 8.03306e-39 + -1.17473e-38 = -3.71422e-39
	(b"10000000011101001100011001010010", b"00000000000000000000000000000000"),
	(b"00000000011110000001101011100110", b"00000000000000110101010010010100"), -- -1.07241e-38 + 1.10299e-38 = 3.05847e-40
	(b"00000000010000000100110001101100", b"00000000000000000000000000000000"),
	(b"10000000010001010011000111001001", b"10000000000001001110010101011101"), -- 5.90489e-39 + -6.35451e-39 = -4.49622e-40
	(b"10000000011111110101101101101100", b"00000000000000000000000000000000"),
	(b"00000000001100010110000000001001", b"10000000010011011111101101100011"), -- -1.16959e-38 + 4.53439e-39 = -7.16151e-39
	(b"10000000000100011101111110100000", b"00000000000000000000000000000000"),
	(b"00000000000001111000110100001000", b"10000000000010100101001010011000"), -- -1.64142e-39 + 6.93441e-40 = -9.47984e-40
	(b"00000000000010101101011000100000", b"00000000000000000000000000000000"),
	(b"10000000010101100101110111100010", b"10000000010010111000011111000010"), -- 9.95169e-40 + -7.93153e-39 = -6.93636e-39
	(b"00000000011000000011100101110110", b"00000000000000000000000000000000"),
	(b"00000000000100011010011001000010", b"00000000011100011101111110111000"), -- 8.83682e-39 + 1.62085e-39 = 1.04577e-38
	(b"00000000001011100010101100000110", b"00000000000000000000000000000000"),
	(b"10000000000101101111010111100101", b"00000000000101110011010100100001"), -- 4.23987e-39 + -2.10859e-39 = 2.13128e-39
	(b"10000000000111001000111100000110", b"00000000000000000000000000000000"),
	(b"00000000000111010001110000000110", b"00000000000000001000110100000000"), -- -2.6227e-39 + 2.67328e-39 = 5.05813e-41
	(b"00000000011011100011101011010011", b"00000000000000000000000000000000"),
	(b"00000000001000000100001010000000", b"00000000100011100111110101010011"), -- 1.0123e-38 + 2.96259e-39 = 1.30856e-38
	(b"00000000011001101000110100100100", b"00000000000000000000000000000000"),
	(b"00000000001001000011011100111010", b"00000000100010101100010001011110"), -- 9.41785e-39 + 3.32589e-39 = 1.27437e-38
	(b"00000000001111011010001000000000", b"00000000000000000000000000000000"),
	(b"00000000001110000101100001100110", b"00000000011101011111101001100110"), -- 5.66008e-39 + 5.1745e-39 = 1.08346e-38
	(b"00000000000101000111100101000000", b"00000000000000000000000000000000"),
	(b"10000000000011101010010000000011", b"00000000000001011101010100111101"), -- 1.88021e-39 + -1.34453e-39 = 5.35673e-40
	(b"00000000011101001100001000001110", b"00000000000000000000000000000000"),
	(b"10000000000000110110011111111101", b"00000000011100010101101000010001"), -- 1.07225e-38 + -3.1281e-40 = 1.04097e-38
	(b"00000000001000010011011011110001", b"00000000000000000000000000000000"),
	(b"10000000001011110110001001111010", b"10000000000011100010101110001001"), -- 3.05028e-39 + -4.3516e-39 = -1.30131e-39
	(b"00000000001100001000011111000110", b"00000000000000000000000000000000"),
	(b"10000000000000101111101011000101", b"00000000001011011000110100000001"), -- 4.45681e-39 + -2.7363e-40 = 4.18318e-39
	(b"10000000000010101001110101001100", b"00000000000000000000000000000000"),
	(b"00000000010110000010100110110101", b"00000000010011011000110001101001"), -- -9.74782e-40 + 8.09649e-39 = 7.1217e-39
	(b"10000000000010110101101011100100", b"00000000000000000000000000000000"),
	(b"00000000011111000101010001111101", b"00000000011100001111100110011001"), -- -1.0428e-39 + 1.14179e-38 = 1.03751e-38
	(b"00000000010001101111010110110000", b"00000000000000000000000000000000"),
	(b"00000000010100000010001010000010", b"00000000100101110001100000110010"), -- 6.51662e-39 + 7.35922e-39 = 1.38758e-38
	(b"00000000000010111100111000111111", b"00000000000000000000000000000000"),
	(b"10000000001000010010111000111110", b"10000000000101010101111111111111"), -- 1.08418e-39 + -3.04716e-39 = -1.96298e-39
	(b"10000000000110000001101001100100", b"00000000000000000000000000000000"),
	(b"10000000011000000011010011010001", b"10000000011110000100111100110101"), -- -2.21352e-39 + -8.83515e-39 = -1.10487e-38
	(b"00000000000010101011010100111011", b"00000000000000000000000000000000"),
	(b"00000000001000011000011000110101", b"00000000001011000011101101110000"), -- 9.83368e-40 + 3.07872e-39 = 4.06208e-39
	(b"00000000010101110000001001100000", b"00000000000000000000000000000000"),
	(b"00000000001000001010101000110001", b"00000000011101111010110010010001"), -- 7.99054e-39 + 2.99979e-39 = 1.09903e-38
	(b"10000000001110010101110101111101", b"00000000000000000000000000000000"),
	(b"00000000000110101110100100101100", b"10000000000111100111010001010001"), -- -5.26816e-39 + 2.47137e-39 = -2.79679e-39
	(b"10000000001001111100110101011010", b"00000000000000000000000000000000"),
	(b"10000000010001000000101110110001", b"10000000011010111101100100001011"), -- -3.65525e-39 + -6.24901e-39 = -9.90426e-39
	(b"00000000011000101011000010010111", b"00000000000000000000000000000000"),
	(b"00000000011000101010101000001010", b"00000000110001010101101010100001"), -- 9.06323e-39 + 9.06088e-39 = 1.81241e-38
	(b"00000000000011010001100100111011", b"00000000000000000000000000000000"),
	(b"00000000010111110000011101111010", b"00000000011011000010000010110101"), -- 1.20291e-39 + 8.72705e-39 = 9.92997e-39
	(b"00000000010000100100100000011111", b"00000000000000000000000000000000"),
	(b"10000000011001110110000010101010", b"10000000001001010001100010001011"), -- 6.08701e-39 + -9.49373e-39 = -3.40672e-39
	(b"10000000000100110011010001000110", b"00000000000000000000000000000000"),
	(b"00000000010010111011001001110101", b"00000000001110000111111000101111"), -- -1.76363e-39 + 6.95168e-39 = 5.18805e-39
	(b"10000000010001010000101010111111", b"00000000000000000000000000000000"),
	(b"10000000001000100010100111000100", b"10000000011001110011010010000011"), -- -6.3405e-39 + -3.13739e-39 = -9.47789e-39
	(b"00000000011001111010001100000111", b"00000000000000000000000000000000"),
	(b"00000000001001110010001100111110", b"00000000100011101100011001000101"), -- 9.51754e-39 + 3.59423e-39 = 1.31118e-38
	(b"10000000010011000011000110011000", b"00000000000000000000000000000000"),
	(b"10000000000100100101000100000110", b"10000000010111101000001010011110"), -- -6.99729e-39 + -1.6821e-39 = -8.67939e-39
	(b"10000000001100001111001011110001", b"00000000000000000000000000000000"),
	(b"10000000010001001011101101100011", b"10000000011101011010111001010100"), -- -4.49525e-39 + -6.31204e-39 = -1.08073e-38
	(b"10000000010011000100111001001010", b"00000000000000000000000000000000"),
	(b"10000000001001100101011101001010", b"10000000011100101010010110010100"), -- -7.00758e-39 + -3.52106e-39 = -1.05286e-38
	(b"10000000001011100001010000111001", b"00000000000000000000000000000000"),
	(b"00000000010110010010000011100111", b"00000000001010110000110010101110"), -- -4.23169e-39 + 8.18516e-39 = 3.95347e-39
	(b"10000000011111110100101101010010", b"00000000000000000000000000000000"),
	(b"00000000001100111011010101010110", b"10000000010010111001010111111100"), -- -1.16901e-38 + 4.74866e-39 = -6.94147e-39
	(b"00000000011100101001111010001101", b"00000000000000000000000000000000"),
	(b"00000000011000100111101111111110", b"00000000110101010001101010001011"), -- 1.05261e-38 + 9.04436e-39 = 1.95705e-38
	(b"00000000001100101001010111110100", b"00000000000000000000000000000000"),
	(b"10000000001010101000111010111011", b"00000000000010000000011100111001"), -- 4.64557e-39 + -3.90829e-39 = 7.37275e-40
	(b"00000000011111000110000010000111", b"00000000000000000000000000000000"),
	(b"10000000000110001010101101100011", b"00000000011000111011010100100100"), -- 1.14222e-38 + -2.26553e-39 = 9.1567e-39
	(b"00000000000100110011101110100101", b"00000000000000000000000000000000"),
	(b"10000000011010100011110111101110", b"10000000010101110000001001001001"), -- 1.76627e-39 + -9.75678e-39 = -7.99051e-39
	(b"00000000010010000110001001100010", b"00000000000000000000000000000000"),
	(b"10000000011110001101011001010101", b"10000000001100000111001111110011"), -- 6.64745e-39 + -1.10971e-38 = -4.4497e-39
	(b"10000000010111010010001000010011", b"00000000000000000000000000000000"),
	(b"00000000001001111101010100001101", b"10000000001101010100110100000110"), -- -8.55292e-39 + 3.65801e-39 = -4.89491e-39
	(b"10000000001111111111110110000111", b"00000000000000000000000000000000"),
	(b"10000000011100011110110011111110", b"10000000101100011110101010000101"), -- -5.87658e-39 + -1.04624e-38 = -1.6339e-38
	(b"10000000010010110111010010110010", b"00000000000000000000000000000000"),
	(b"10000000010000100101010010110101", b"10000000100011011100100101100111"), -- -6.92952e-39 + -6.09153e-39 = -1.30211e-38
	(b"00000000001011011000101111010100", b"00000000000000000000000000000000"),
	(b"10000000000100100100010011000110", b"00000000000110110100011100001110"), -- 4.18276e-39 + -1.67771e-39 = 2.50505e-39
	(b"10000000000111001000010010110111", b"00000000000000000000000000000000"),
	(b"00000000000111010100111101111011", b"00000000000000001100101011000100"), -- -2.619e-39 + 2.69174e-39 = 7.27386e-41
	(b"10000000011001110101101101001011", b"00000000000000000000000000000000"),
	(b"10000000001111011010110101001010", b"10000000101001010000100010010101"), -- -9.49181e-39 + -5.66413e-39 = -1.51559e-38
	(b"10000000001110011110011000011000", b"00000000000000000000000000000000"),
	(b"00000000001110010000010101110010", b"10000000000000001110000010100110"), -- -5.31717e-39 + 5.23658e-39 = -8.05887e-41
	(b"10000000001010110000110110010000", b"00000000000000000000000000000000"),
	(b"10000000001100110010010011011111", b"10000000010111100011001001101111"), -- -3.95379e-39 + -4.69684e-39 = -8.65063e-39
	(b"00000000011010100101011010101110", b"00000000000000000000000000000000"),
	(b"00000000001011101100010000000010", b"00000000100110010001101010110000"), -- 9.76566e-39 + 4.29475e-39 = 1.40604e-38
	(b"00000000011100111000110001110001", b"00000000000000000000000000000000"),
	(b"00000000000111110000001100001010", b"00000000100100101000111101111011"), -- 1.06115e-38 + 2.84799e-39 = 1.34595e-38
	(b"00000000001111100111000010101011", b"00000000000000000000000000000000"),
	(b"00000000000011100101010101100111", b"00000000010011001100011000010010"), -- 5.73422e-39 + 1.31633e-39 = 7.05055e-39
	(b"00000000000110000011101010110001", b"00000000000000000000000000000000"),
	(b"00000000001000111000011010011010", b"00000000001110111100000101001011"), -- 2.22511e-39 + 3.26253e-39 = 5.48763e-39
	(b"00000000001000110100111011001000", b"00000000000000000000000000000000"),
	(b"00000000011110100001101111010110", b"00000000100111010110101010011110"), -- 3.2425e-39 + 1.12139e-38 = 1.44564e-38
	(b"00000000000100111010011000100010", b"00000000000000000000000000000000"),
	(b"10000000001001010100111010110000", b"10000000000100011010100010001110"), -- 1.80447e-39 + -3.42614e-39 = -1.62167e-39
	(b"00000000011010001011111100100001", b"00000000000000000000000000000000"),
	(b"10000000001101011101010100000101", b"00000000001100101110101000011100"), -- 9.61946e-39 + -4.9437e-39 = 4.67576e-39
	(b"00000000011001001101010000010001", b"00000000000000000000000000000000"),
	(b"00000000011011000000010110111100", b"00000000110100001101100111001101"), -- 9.25962e-39 + 9.92029e-39 = 1.91799e-38
	(b"10000000000101001101101010000001", b"00000000000000000000000000000000"),
	(b"10000000001100101111001011100001", b"10000000010001111100110101100010"), -- -1.91509e-39 + -4.6789e-39 = -6.594e-39
	(b"00000000000111010011011101110100", b"00000000000000000000000000000000"),
	(b"10000000001111001001010111110010", b"10000000000111110101111001111110"), -- 2.68312e-39 + -5.56392e-39 = -2.8808e-39
	(b"00000000000000111111010101111101", b"00000000000000000000000000000000"),
	(b"10000000010110001000000101011100", b"10000000010101001000101111011111"), -- 3.63571e-40 + -8.12793e-39 = -7.76436e-39
	(b"10000000000011000100010010110110", b"00000000000000000000000000000000"),
	(b"00000000001101011110110010001000", b"00000000001010011010011111010010"), -- -1.12667e-39 + 4.95213e-39 = 3.82546e-39
	(b"10000000010111110010100000110000", b"00000000000000000000000000000000"),
	(b"00000000011001000001000010001111", b"00000000000001001110100001011111"), -- -8.73879e-39 + 9.18949e-39 = 4.50701e-40
	(b"00000000001011010110101010110010", b"00000000000000000000000000000000"),
	(b"00000000000001001100100011100111", b"00000000001100100011001110011001"), -- 4.17087e-39 + 4.39412e-40 = 4.61028e-39
	(b"10000000011000110111111100110111", b"00000000000000000000000000000000"),
	(b"10000000001100011110101001001010", b"10000000100101010110100110000001"), -- -9.13735e-39 + -4.58399e-39 = -1.37213e-38
	(b"10000000011101111111101110110101", b"00000000000000000000000000000000"),
	(b"10000000011100111101110111100011", b"10000000111010111101100110011000"), -- -1.10187e-38 + -1.06407e-38 = -2.16594e-38
	(b"00000000011100001000011010100000", b"00000000000000000000000000000000"),
	(b"00000000011111110111001100001110", b"00000000111011111111100110101110"), -- 1.03339e-38 + 1.17044e-38 = 2.20383e-38
	(b"00000000000101010000101100110111", b"00000000000000000000000000000000"),
	(b"10000000001011101001011000111001", b"10000000000110011000101100000010"), -- 1.93257e-39 + -4.27832e-39 = -2.34575e-39
	(b"00000000001100001111110001100111", b"00000000000000000000000000000000"),
	(b"10000000011110100001001000000001", b"10000000010010010001010110011010"), -- 4.49865e-39 + -1.12104e-38 = -6.71174e-39
	(b"10000000010101100000010011011011", b"00000000000000000000000000000000"),
	(b"00000000000011000011010110101100", b"10000000010010011100111100101111"), -- -7.89959e-39 + 1.12128e-39 = -6.77831e-39
	(b"10000000001000101111100101100011", b"00000000000000000000000000000000"),
	(b"10000000010101110000100110111101", b"10000000011110100000001100100000"), -- -3.21187e-39 + -7.99318e-39 = -1.12051e-38
	(b"10000000001111001011011000110011", b"00000000000000000000000000000000"),
	(b"10000000000100101110100011001011", b"10000000010011111001111011111110"), -- -5.57549e-39 + -1.73655e-39 = -7.31204e-39
	(b"10000000011011010011000100110000", b"00000000000000000000000000000000"),
	(b"10000000010001001011110111011001", b"10000000101100011110111100001001"), -- -1.00277e-38 + -6.31292e-39 = -1.63406e-38
	(b"10000000000111011000001110110110", b"00000000000000000000000000000000"),
	(b"00000000011100110011100011000111", b"00000000010101011011010100010001"), -- -2.71048e-39 + 1.05814e-38 = 7.87097e-39
	(b"10000000011010000100010100010000", b"00000000000000000000000000000000"),
	(b"10000000010110101110101000000000", b"10000000110000110010111100010000"), -- -9.57567e-39 + -8.34914e-39 = -1.79248e-38
	(b"10000000001010011000111010111011", b"00000000000000000000000000000000"),
	(b"10000000001000000111101100110001", b"10000000010010100000100111101100"), -- -3.81646e-39 + -2.98293e-39 = -6.79939e-39
	(b"10000000000010111000010000100110", b"00000000000000000000000000000000"),
	(b"10000000011110000011011111111000", b"10000000100000111011110000011110"), -- -1.0576e-39 + -1.10403e-38 = -1.20979e-38
	(b"00000000011110001100101100001101", b"00000000000000000000000000000000"),
	(b"10000000010101111010111001010010", b"00000000001000010001110010111011"), -- 1.10931e-38 + -8.05222e-39 = 3.04088e-39
	(b"10000000000011100010010101000000", b"00000000000000000000000000000000"),
	(b"00000000001110111011010000111101", b"00000000001011011000111011111101"), -- -1.29906e-39 + 5.48295e-39 = 4.18389e-39
	(b"10000000001111100101101111101000", b"00000000000000000000000000000000"),
	(b"00000000001101011011101010001011", b"10000000000010001010000101011101"), -- -5.72677e-39 + 4.9342e-39 = -7.9257e-40
	(b"00000000011111110111111111110110", b"00000000000000000000000000000000"),
	(b"00000000011100010001110101110111", b"00000000111100001001110101101101"), -- 1.1709e-38 + 1.0388e-38 = 2.2097e-38
	(b"00000000010010111010100010010000", b"00000000000000000000000000000000"),
	(b"00000000010110010011101111111011", b"00000000101001001110010010001011"), -- 6.94813e-39 + 8.19488e-39 = 1.5143e-38
	(b"10000000000010000011001100100000", b"00000000000000000000000000000000"),
	(b"10000000000100001110011100000010", b"10000000000110010001101000100010"), -- -7.53024e-40 + -1.55224e-39 = -2.30526e-39
	(b"10000000000111001000111110111111", b"00000000000000000000000000000000"),
	(b"10000000010000100100110010001111", b"10000000010111101101110001001110"), -- -2.62296e-39 + -6.08861e-39 = -8.71157e-39
	(b"10000000001111001110000100010011", b"00000000000000000000000000000000"),
	(b"00000000001100101010010010100000", b"10000000000010100011110001110011"), -- -5.59087e-39 + 4.65083e-39 = -9.4004e-40
	(b"00000000011000110110000111100000", b"00000000000000000000000000000000"),
	(b"00000000011111100100111011000010", b"00000000111000011011000010100010"), -- 9.12683e-39 + 1.15995e-38 = 2.07264e-38
	(b"10000000010010101000010110000010", b"00000000000000000000000000000000"),
	(b"10000000010001101001100100010100", b"10000000100100010001111010010110"), -- -6.84372e-39 + -6.4834e-39 = -1.33271e-38
	(b"10000000011111101100101011011000", b"00000000000000000000000000000000"),
	(b"00000000000111010101001100011101", b"10000000011000010111011110111011"), -- -1.1644e-38 + 2.69304e-39 = -8.95099e-39
	(b"00000000011011001000011101101001", b"00000000000000000000000000000000"),
	(b"00000000011101101100110101000001", b"00000000111000110101010010101010"), -- 9.96681e-39 + 1.09102e-38 = 2.0877e-38
	(b"00000000000001110111000110110010", b"00000000000000000000000000000000"),
	(b"10000000001100000101011101010011", b"10000000001010001110010110100001"), -- 6.83635e-40 + -4.43943e-39 = -3.7558e-39
	(b"10000000000010110100001100000010", b"00000000000000000000000000000000"),
	(b"00000000001101111101010010111010", b"00000000001011001001000110111000"), -- -1.03423e-39 + 5.12726e-39 = 4.09304e-39
	(b"10000000010000001100011011101000", b"00000000000000000000000000000000"),
	(b"00000000011100101110110110111001", b"00000000001100100010011011010001"), -- -5.94883e-39 + 1.05545e-38 = 4.6057e-39
	(b"00000000011111001000110001010101", b"00000000000000000000000000000000"),
	(b"10000000001101100110100011000010", b"00000000010001100010001110010011"), -- 1.14379e-38 + -4.9967e-39 = 6.44125e-39
	(b"10000000010001100010111010100001", b"00000000000000000000000000000000"),
	(b"10000000010110000100010101010000", b"10000000100111100111001111110001"), -- -6.44521e-39 + -8.10639e-39 = -1.45516e-38
	(b"00000000010010100001100110001010", b"00000000000000000000000000000000"),
	(b"00000000000101000111000110000000", b"00000000010111101000101100001010"), -- 6.80499e-39 + 1.87743e-39 = 8.68241e-39
	(b"10000000000111101101111110101100", b"00000000000000000000000000000000"),
	(b"00000000010111100011001010010010", b"00000000001111110101001011100110"), -- -2.8353e-39 + 8.65068e-39 = 5.81537e-39
	(b"00000000000000111011101101100011", b"00000000000000000000000000000000"),
	(b"10000000001000001101010101011011", b"10000000000111010001100111111000"), -- 3.42728e-40 + -3.01527e-39 = -2.67255e-39
	(b"10000000010011001101100000100100", b"00000000000000000000000000000000"),
	(b"10000000010101110100010111011110", b"10000000101001000001111000000010"), -- -7.05703e-39 + -8.01475e-39 = -1.50718e-38
	(b"00000000000000110000011101101111", b"00000000000000000000000000000000"),
	(b"00000000001000001011000000001111", b"00000000001000111011011101111110"), -- 2.78173e-40 + 3.00189e-39 = 3.28007e-39
	(b"00000000001111100000101101111011", b"00000000000000000000000000000000"),
	(b"10000000001001010110000000111011", b"00000000000110001010101101000000"), -- 5.69792e-39 + -3.43243e-39 = 2.26548e-39
	(b"10000000001101110010100101011100", b"00000000000000000000000000000000"),
	(b"00000000001010001111101000100100", b"10000000000011100010111100111000"), -- -5.06579e-39 + 3.76315e-39 = -1.30264e-39
	(b"00000000000110111011100110100101", b"00000000000000000000000000000000"),
	(b"10000000000000010101011101111111", b"00000000000110100110001000100110"), -- 2.54616e-39 + -1.23223e-40 = 2.42293e-39
	(b"00000000001001001111010110011100", b"00000000000000000000000000000000"),
	(b"10000000001000001000111000100100", b"00000000000001000110011101111000"), -- 3.39419e-39 + -2.98973e-39 = 4.0446e-40
	(b"10000000001010110100101111011111", b"00000000000000000000000000000000"),
	(b"10000000000011111001100010101100", b"10000000001110101110010010001011"), -- -3.97614e-39 + -1.4323e-39 = -5.40844e-39
	(b"10000000001110110000101001100010", b"00000000000000000000000000000000"),
	(b"10000000000010011001101010101101", b"10000000010001001010010100001111"), -- -5.42202e-39 + -8.82007e-40 = -6.30403e-39
	(b"10000000001001110000000101100110", b"00000000000000000000000000000000"),
	(b"10000000001011101110011000011001", b"10000000010101011110011101111111"), -- -3.58209e-39 + -4.30698e-39 = -7.88906e-39
	(b"00000000010011000010100101001010", b"00000000000000000000000000000000"),
	(b"10000000011001110000111011010000", b"10000000000110101110010110000110"), -- 6.99431e-39 + -9.46437e-39 = -2.47006e-39
	(b"00000000000110000011111010101010", b"00000000000000000000000000000000"),
	(b"10000000011100011101110110000011", b"10000000010110011001111011011001"), -- 2.22653e-39 + -1.04569e-38 = -8.23034e-39
	(b"10000000001101110011010111001010", b"00000000000000000000000000000000"),
	(b"00000000001100111111100011001001", b"10000000000000110011110100000001"), -- -5.07025e-39 + 4.77286e-39 = -2.97391e-40
	(b"10000000011111001101110010110110", b"00000000000000000000000000000000"),
	(b"00000000000000101110111001011010", b"10000000011110011110111001011100"), -- -1.14668e-38 + 2.69175e-40 = -1.11976e-38
	(b"00000000011111010101110001110000", b"00000000000000000000000000000000"),
	(b"10000000011001100010101100011111", b"00000000000101110011000101010001"), -- 1.15126e-38 + -9.38269e-39 = 2.12991e-39
	(b"10000000010001000101110010011010", b"00000000000000000000000000000000"),
	(b"00000000000001100010111110011101", b"10000000001111100010110011111101"), -- -6.27803e-39 + 5.68093e-40 = -5.70994e-39
	(b"00000000000101011100011001111101", b"00000000000000000000000000000000"),
	(b"00000000000101011100111011010001", b"00000000001010111001010101001110"), -- 1.99975e-39 + 2.00274e-39 = 4.00249e-39
	(b"10000000001001011000001011000001", b"00000000000000000000000000000000"),
	(b"00000000010011010001000110111100", b"00000000001001111000111011111011"), -- -3.44482e-39 + 7.0777e-39 = 3.63288e-39
	(b"10000000001111100001111011101100", b"00000000000000000000000000000000"),
	(b"00000000000111001100001100110101", b"10000000001000010101101110110111"), -- -5.70489e-39 + 2.64142e-39 = -3.06347e-39
	(b"10000000001101011000111111010101", b"00000000000000000000000000000000"),
	(b"00000000001011100001001110001111", b"10000000000001110111110001000110"), -- -4.91888e-39 + 4.23145e-39 = -6.87429e-40
	(b"10000000001001001001110011100100", b"00000000000000000000000000000000"),
	(b"10000000011101110000011101011000", b"10000000100110111010010000111100"), -- -3.36236e-39 + -1.09311e-38 = -1.42934e-38
	(b"00000000011110001000010010111100", b"00000000000000000000000000000000"),
	(b"00000000000011100011101011110100", b"00000000100001101011111110110000"), -- 1.10679e-38 + 1.30685e-39 = 1.23747e-38
	(b"10000000000000101101101100001000", b"00000000000000000000000000000000"),
	(b"10000000011110101100110001110001", b"10000000011111011010011101111001"), -- -2.62245e-40 + -1.12773e-38 = -1.15395e-38
	(b"10000000011000110101011001001011", b"00000000000000000000000000000000"),
	(b"10000000011001101011001011111001", b"10000000110010100000100101000100"), -- -9.12267e-39 + -9.43142e-39 = -1.85541e-38
	(b"10000000010101000001000011110110", b"00000000000000000000000000000000"),
	(b"10000000000011011101101001011001", b"10000000011000011110101101001111"), -- -7.72027e-39 + -1.27219e-39 = -8.99246e-39
	(b"00000000001010000011100011000101", b"00000000000000000000000000000000"),
	(b"00000000000001101011010000100010", b"00000000001011101110110011100111"), -- 3.69378e-39 + 6.15632e-40 = 4.30942e-39
	(b"10000000000001011010000101001010", b"00000000000000000000000000000000"),
	(b"10000000000000011010010110101101", b"10000000000001110100011011110111"), -- -5.17037e-40 + -1.51269e-40 = -6.68306e-40
	(b"10000000001001000011010000001010", b"00000000000000000000000000000000"),
	(b"00000000000011101111001111001001", b"10000000000101010100000001000001"), -- -3.32475e-39 + 1.37315e-39 = -1.9516e-39
	(b"10000000001011101000110101100001", b"00000000000000000000000000000000"),
	(b"00000000011010011011010010101011", b"00000000001110110010011101001010"), -- -4.27515e-39 + 9.70754e-39 = 5.43239e-39
	(b"10000000000110011101001001001011", b"00000000000000000000000000000000"),
	(b"10000000010001011100111111101110", b"10000000010111111010001000111001"), -- -2.37133e-39 + -6.41124e-39 = -8.78257e-39
	(b"00000000000011000000110011100101", b"00000000000000000000000000000000"),
	(b"00000000000011100001010111001101", b"00000000000110100010001010110010"), -- 1.10665e-39 + 1.29352e-39 = 2.40017e-39
	(b"10000000000101011110011010110111", b"00000000000000000000000000000000"),
	(b"00000000011000011011110001010000", b"00000000010010111101010110011001"), -- -2.01131e-39 + 8.9756e-39 = 6.96429e-39
	(b"00000000000000001010001011111001", b"00000000000000000000000000000000"),
	(b"10000000000011001101010011001111", b"10000000000011000011000111010110"), -- 5.84636e-41 + -1.17837e-39 = -1.1199e-39
	(b"00000000001110001000001110101000", b"00000000000000000000000000000000"),
	(b"00000000010001111100011111011111", b"00000000100000000100101110000111"), -- 5.19002e-39 + 6.59202e-39 = 1.1782e-38
	(b"10000000000001101110110100001000", b"00000000000000000000000000000000"),
	(b"00000000011011000000010100011011", b"00000000011001010001100000010011"), -- -6.36044e-40 + 9.92007e-39 = 9.28402e-39
	(b"00000000011001101100001000000001", b"00000000000000000000000000000000"),
	(b"00000000011110001010011010000111", b"00000000110111110110100010001000"), -- 9.43682e-39 + 1.108e-38 = 2.05168e-38
	(b"10000000010000010100000001010110", b"00000000000000000000000000000000"),
	(b"00000000001111011011000111001000", b"10000000000000111000111010001110"), -- -5.99239e-39 + 5.66574e-39 = -3.26645e-40
	(b"10000000000111010101000001101111", b"00000000000000000000000000000000"),
	(b"10000000011100111000000111010010", b"10000000100100001101001001000001"), -- -2.69208e-39 + -1.06077e-38 = -1.32997e-38
	(b"10000000000000001101010100010100", b"00000000000000000000000000000000"),
	(b"10000000011010000111011110100110", b"10000000011010010100110010111010"), -- -7.6438e-41 + -9.59381e-39 = -9.67025e-39
	(b"10000000011000110010110110100001", b"00000000000000000000000000000000"),
	(b"00000000011010001001101100111010", b"00000000000001010110110110011001"), -- -9.10808e-39 + 9.60658e-39 = 4.98494e-40
	(b"00000000011011000110011010110001", b"00000000000000000000000000000000"),
	(b"10000000011110111000110011110110", b"10000000000011110010011001000101"), -- 9.95507e-39 + -1.13463e-38 = -1.39126e-39
	(b"00000000011000000011000001000010", b"00000000000000000000000000000000"),
	(b"00000000011011100101000010001110", b"00000000110011101000000011010000"), -- 8.83352e-39 + 1.01308e-38 = 1.89643e-38
	(b"00000000001001011001011011110110", b"00000000000000000000000000000000"),
	(b"00000000010010100000110100001101", b"00000000011011111010010000000011"), -- 3.45207e-39 + 6.80051e-39 = 1.02526e-38
	(b"10000000011010001101011011100010", b"00000000000000000000000000000000"),
	(b"00000000011101010111011010011110", b"00000000000011001001111110111100"), -- -9.62798e-39 + 1.07873e-38 = 1.15933e-39
	(b"00000000001111001000111111011111", b"00000000000000000000000000000000"),
	(b"00000000011100100110001100111110", b"00000000101011101111001100011101"), -- 5.56174e-39 + 1.05048e-38 = 1.60666e-38
	(b"00000000001001010010011111111011", b"00000000000000000000000000000000"),
	(b"10000000000100000001111100110001", b"00000000000101010000100011001010"), -- 3.41226e-39 + -1.48056e-39 = 1.9317e-39
	(b"10000000010110001001001100000101", b"00000000000000000000000000000000"),
	(b"00000000001010101001011001110100", b"10000000001011011111110010010001"), -- -8.13426e-39 + 3.91106e-39 = -4.2232e-39
	(b"10000000001010110111000101001101", b"00000000000000000000000000000000"),
	(b"10000000010110010000101110101111", b"10000000100001000111110011111100"), -- -3.98957e-39 + -8.17755e-39 = -1.21671e-38
	(b"10000000001011100111110111111010", b"00000000000000000000000000000000"),
	(b"00000000000000110111011111111001", b"10000000001010110000011000000001"), -- -4.26962e-39 + 3.18545e-40 = -3.95108e-39
	(b"10000000001100100011110101011000", b"00000000000000000000000000000000"),
	(b"10000000001000011010100000100100", b"10000000010100111110010101111100"), -- -4.61378e-39 + -3.09089e-39 = -7.70467e-39
	(b"10000000001001100111011111101110", b"00000000000000000000000000000000"),
	(b"00000000011100000101100000100010", b"00000000010010011110000000110100"), -- -3.53277e-39 + 1.03172e-38 = 6.78442e-39
	(b"10000000000100110011011011110101", b"00000000000000000000000000000000"),
	(b"00000000010001010000100111011001", b"00000000001100011101001011100100"), -- -1.76459e-39 + 6.34018e-39 = 4.57559e-39
	(b"10000000010010010110100011011101", b"00000000000000000000000000000000"),
	(b"00000000001101000100101010000110", b"10000000000101010001111001010111"), -- -6.74161e-39 + 4.80218e-39 = -1.93943e-39
	(b"10000000001011101101101000010011", b"00000000000000000000000000000000"),
	(b"00000000011001000111111101000111", b"00000000001101011010010100110100"), -- -4.30266e-39 + 9.22921e-39 = 4.92655e-39
	(b"10000000001100010001010100010101", b"00000000000000000000000000000000"),
	(b"10000000010110111100100101010110", b"10000000100011001101111001101011"), -- -4.5075e-39 + -8.42926e-39 = -1.29368e-38
	(b"10000000000100011011111110100000", b"00000000000000000000000000000000"),
	(b"00000000001100000011100100111111", b"00000000000111100111100110011111"), -- -1.62995e-39 + 4.42864e-39 = 2.79869e-39
	(b"10000000011111101100110000101011", b"00000000000000000000000000000000"),
	(b"00000000000110110110111101000101", b"10000000011000110101110011100110"), -- -1.16445e-38 + 2.51947e-39 = -9.12504e-39
	(b"00000000010110101110100001111001", b"00000000000000000000000000000000"),
	(b"10000000000011101000101010001100", b"00000000010011000101110111101101"), -- 8.34859e-39 + -1.3354e-39 = 7.01319e-39
	(b"00000000000010001010010011110000", b"00000000000000000000000000000000"),
	(b"10000000000110011011010101001011", b"10000000000100010001000001011011"), -- 7.93852e-40 + -2.36092e-39 = -1.56707e-39
	(b"10000000000110001101101100101111", b"00000000000000000000000000000000"),
	(b"00000000001101001001001111100000", b"00000000000110111011100010110001"), -- -2.28268e-39 + 4.82849e-39 = 2.54581e-39
	(b"00000000001010001000110110010101", b"00000000000000000000000000000000"),
	(b"10000000001110101000000010110100", b"10000000000100011111001100011111"), -- 3.72421e-39 + -5.37263e-39 = -1.64842e-39
	(b"00000000010011100100101111001001", b"00000000000000000000000000000000"),
	(b"00000000001110101101101111011011", b"00000000100010010010011110100100"), -- 7.19036e-39 + 5.40533e-39 = 1.25957e-38
	(b"10000000000000100010101111111111", b"00000000000000000000000000000000"),
	(b"00000000001000101100100111010100", b"00000000001000001001110111010101"), -- -1.99454e-40 + 3.19481e-39 = 2.99536e-39
	(b"00000000010000101111111001011101", b"00000000000000000000000000000000"),
	(b"10000000010011100001111001101101", b"10000000000010110010000000010000"), -- 6.15239e-39 + -7.17408e-39 = -1.02169e-39
	(b"10000000011010010011000111001110", b"00000000000000000000000000000000"),
	(b"10000000000110100011100010010011", b"10000000100000110110101001100001"), -- -9.66059e-39 + -2.40802e-39 = -1.20686e-38
	(b"10000000010010111101110110000101", b"00000000000000000000000000000000"),
	(b"00000000011000110101010110101001", b"00000000000101110111100000100100"), -- -6.96713e-39 + 9.12244e-39 = 2.15531e-39
	(b"00000000010100101011110011111101", b"00000000000000000000000000000000"),
	(b"10000000011000011001001100100100", b"10000000000011101101011000100111"), -- 7.59831e-39 + -8.96083e-39 = -1.36252e-39
	(b"00000000011111011001001101100101", b"00000000000000000000000000000000"),
	(b"10000000010111010100001110110110", b"00000000001000000100111110101111"), -- 1.15323e-38 + -8.56499e-39 = 2.96732e-39
	(b"00000000001000110000110011100111", b"00000000000000000000000000000000"),
	(b"10000000010000001101000110101100", b"10000000000111011100010011000101"), -- 3.21887e-39 + -5.95269e-39 = -2.73382e-39
	(b"10000000010111010111011010011001", b"00000000000000000000000000000000"),
	(b"10000000010001101110101111011110", b"10000000101001000110001001110111"), -- -8.58325e-39 + -6.5131e-39 = -1.50963e-38
	(b"10000000001010110101111100110110", b"00000000000000000000000000000000"),
	(b"00000000001011100110001100011011", b"00000000000000110000001111100101"), -- -3.98308e-39 + 4.25999e-39 = 2.76904e-40
	(b"00000000000101001100000111110111", b"00000000000000000000000000000000"),
	(b"00000000010111011100001110110010", b"00000000011100101000010110101001"), -- 1.90629e-39 + 8.6109e-39 = 1.05172e-38
	(b"00000000011011001110101101110110", b"00000000000000000000000000000000"),
	(b"10000000011101101101001010011111", b"10000000000010011110011100101001"), -- 1.00027e-38 + -1.09121e-38 = -9.09444e-40
	(b"00000000011101000011111100100001", b"00000000000000000000000000000000"),
	(b"00000000010000001001111111000010", b"00000000101101001101111011100011"), -- 1.06756e-38 + 5.93478e-39 = 1.66103e-38
	(b"10000000001100000000101010001010", b"00000000000000000000000000000000"),
	(b"10000000011111010100100000010011", b"10000000101011010101001010011101"), -- -4.41188e-39 + -1.15053e-38 = -1.59172e-38
	(b"10000000000010000010000010101101", b"00000000000000000000000000000000"),
	(b"10000000001111001111110000001011", b"10000000010001010001110010111000"), -- -7.46406e-40 + -5.60055e-39 = -6.34695e-39
	(b"00000000000101000111101010100011", b"00000000000000000000000000000000"),
	(b"00000000010111111000010000011100", b"00000000011100111111111010111111"), -- 1.8807e-39 + 8.77176e-39 = 1.06525e-38
	(b"10000000011010111100010101001110", b"00000000000000000000000000000000"),
	(b"00000000011110011111110110111000", b"00000000000011100011100001101010"), -- -9.89718e-39 + 1.12031e-38 = 1.30593e-39
	(b"00000000011000100000001101111011", b"00000000000000000000000000000000"),
	(b"00000000011011101100101110011000", b"00000000110100001100111100010011"), -- 9.00113e-39 + 1.01749e-38 = 1.91761e-38
	(b"00000000001101100111101011000101", b"00000000000000000000000000000000"),
	(b"10000000010001000010010100010100", b"10000000000011011010101001001111"), -- 5.00316e-39 + -6.25811e-39 = -1.25496e-39
	(b"00000000010010011111000110011001", b"00000000000000000000000000000000"),
	(b"00000000001010110011011001010000", b"00000000011101010010011111101001"), -- 6.79066e-39 + 3.96841e-39 = 1.07591e-38
	(b"10000000010100000001110011000001", b"00000000000000000000000000000000"),
	(b"00000000010101010000011011100010", b"00000000000001001110101000100001"), -- -7.35715e-39 + 7.80849e-39 = 4.51332e-40
	(b"10000000011110011110000101001110", b"00000000000000000000000000000000"),
	(b"00000000000101101111000101001001", b"10000000011000101111000000000101"), -- -1.11929e-38 + 2.10694e-39 = -9.08598e-39
	(b"00000000001000101101101011111101", b"00000000000000000000000000000000"),
	(b"00000000010000011001010100011101", b"00000000011001000111000000011010"), -- 3.20097e-39 + 6.0228e-39 = 9.22376e-39
	(b"10000000001100000010111010100011", b"00000000000000000000000000000000"),
	(b"10000000001000101010111110010011", b"10000000010100101101111000110110"), -- -4.42483e-39 + -3.18539e-39 = -7.61022e-39
	(b"00000000011010000001000000101100", b"00000000000000000000000000000000"),
	(b"10000000010001011111101000001001", b"00000000001000100001011000100011"), -- 9.55669e-39 + -6.42634e-39 = 3.13035e-39
	(b"10000000001101111011000001010010", b"00000000000000000000000000000000"),
	(b"00000000000111001000011111101100", b"10000000000110110010100001100110"), -- -5.1142e-39 + 2.62015e-39 = -2.49405e-39
	(b"00000000011011110000000101110011", b"00000000000000000000000000000000"),
	(b"10000000011011001001110100100000", b"00000000000000100110010001010011"), -- 1.01943e-38 + -9.9746e-39 = 2.19661e-40
	(b"00000000000111111011011110011111", b"00000000000000000000000000000000"),
	(b"00000000011001010001010111111000", b"00000000100001001100110110010111"), -- 2.91277e-39 + 9.28327e-39 = 1.2196e-38
	(b"00000000010110001101111100010000", b"00000000000000000000000000000000"),
	(b"00000000010001101010110011010010", b"00000000100111111000101111100010"), -- 8.16154e-39 + 6.49048e-39 = 1.4652e-38
	(b"10000000001000100110100101001001", b"00000000000000000000000000000000"),
	(b"00000000010111100100000111100101", b"00000000001110111101100010011100"), -- -3.16018e-39 + 8.65618e-39 = 5.496e-39
	(b"00000000000011011001111101101111", b"00000000000000000000000000000000"),
	(b"10000000011011100011001000000001", b"10000000011000001001001010010010"), -- 1.25106e-39 + -1.01198e-38 = -8.86879e-39
	(b"00000000011100001100001100010010", b"00000000000000000000000000000000"),
	(b"10000000001011000001001101011011", b"00000000010001001010111110110111"), -- 1.03556e-38 + -4.04771e-39 = 6.30785e-39
	(b"10000000010110011111011011010011", b"00000000000000000000000000000000"),
	(b"00000000011110000000001000001001", b"00000000000111100000101100110110"), -- -8.2619e-39 + 1.1021e-38 = 2.75909e-39
	(b"10000000001010110101000111000001", b"00000000000000000000000000000000"),
	(b"10000000011110011011110011001111", b"10000000101001010000111010010000"), -- -3.97825e-39 + -1.11798e-38 = -1.51581e-38
	(b"00000000011010110010001010101110", b"00000000000000000000000000000000"),
	(b"00000000000001101011111010101100", b"00000000011100011110000101011010"), -- 9.83884e-39 + 6.19413e-40 = 1.04583e-38
	(b"00000000010011000100010101000010", b"00000000000000000000000000000000"),
	(b"00000000011001100111001110001101", b"00000000101100101011100011001111"), -- 7.00434e-39 + 9.40867e-39 = 1.6413e-38
	(b"00000000010011011100101010101100", b"00000000000000000000000000000000"),
	(b"10000000000011011111100100010100", b"00000000001111111101000110011000"), -- 7.14404e-39 + -1.28321e-39 = 5.86082e-39
	(b"10000000011100001000101111100000", b"00000000000000000000000000000000"),
	(b"00000000000111000111010001101011", b"10000000010101000001011101110101"), -- -1.03358e-38 + 2.61316e-39 = -7.7226e-39
	(b"10000000011110001011010011001001", b"00000000000000000000000000000000"),
	(b"10000000001010001010111111111100", b"10000000101000010110010011000101"), -- -1.10851e-38 + -3.73655e-39 = -1.48217e-38
	(b"10000000010111101011110101100001", b"00000000000000000000000000000000"),
	(b"00000000001000100100011100010110", b"10000000001111000111011001001011"), -- -8.70047e-39 + 3.14791e-39 = -5.55257e-39
	(b"00000000010011001101101100011100", b"00000000000000000000000000000000"),
	(b"10000000000101101010101101100101", b"00000000001101100010111110110111"), -- 7.0581e-39 + -2.08187e-39 = 4.97623e-39
	(b"00000000010001010101111100011010", b"00000000000000000000000000000000"),
	(b"10000000010100100110101101111000", b"10000000000011010000110001011110"), -- 6.37077e-39 + -7.56906e-39 = -1.1983e-39
	(b"00000000001111001110111011001011", b"00000000000000000000000000000000"),
	(b"00000000011001001110101110011001", b"00000000101000011101101001100100"), -- 5.59579e-39 + 9.26807e-39 = 1.48639e-38
	(b"00000000001100100100001001001100", b"00000000000000000000000000000000"),
	(b"00000000001100101011110011010100", b"00000000011001001111111100100000"), -- 4.61556e-39 + 4.65951e-39 = 9.27507e-39
	(b"10000000010110100010010010011010", b"00000000000000000000000000000000"),
	(b"00000000011111010011010110001000", b"00000000001000110001000011101110"), -- -8.27832e-39 + 1.14986e-38 = 3.22032e-39
	(b"10000000000111100101100011000001", b"00000000000000000000000000000000"),
	(b"00000000010010000010010110110010", b"00000000001010011100110011110001"), -- -2.7869e-39 + 6.62568e-39 = 3.83877e-39
	(b"00000000011000010010000100001100", b"00000000000000000000000000000000"),
	(b"00000000001100101001101011011100", b"00000000100100111011101111101000"), -- 8.9199e-39 + 4.64733e-39 = 1.35672e-38
	(b"00000000000010111011000001110000", b"00000000000000000000000000000000"),
	(b"10000000001111110000001111010101", b"10000000001100110101001101100101"), -- 1.07348e-39 + -5.78701e-39 = -4.71353e-39
	(b"00000000011101010000000011101011", b"00000000000000000000000000000000"),
	(b"10000000010111111010001100001001", b"00000000000101010101110111100010"), -- 1.07451e-38 + -8.78286e-39 = 1.96222e-39
	(b"10000000000011001111001100000110", b"00000000000000000000000000000000"),
	(b"00000000001110000010100101111111", b"00000000001010110011011001111001"), -- -1.18921e-39 + 5.15767e-39 = 3.96847e-39
	(b"00000000011001100110011010000110", b"00000000000000000000000000000000"),
	(b"00000000011010010101110001110110", b"00000000110011111100001011111100"), -- 9.404e-39 + 9.6759e-39 = 1.90799e-38
	(b"10000000010110101000011011000101", b"00000000000000000000000000000000"),
	(b"00000000000100110110110011111001", b"10000000010001110001100111001100"), -- -8.31354e-39 + 1.78397e-39 = -6.52957e-39
	(b"10000000011001101110110101000010", b"00000000000000000000000000000000"),
	(b"10000000001010111001100101101101", b"10000000100100101000011010101111"), -- -9.45233e-39 + -4.00397e-39 = -1.34563e-38
	(b"10000000010100011001111110001010", b"00000000000000000000000000000000"),
	(b"10000000000001100100100011110000", b"10000000010101111110100001111010"), -- -7.49591e-39 + -5.77178e-40 = -8.07309e-39
	(b"10000000010001111100111000101010", b"00000000000000000000000000000000"),
	(b"10000000010011101010110010101110", b"10000000100101100111101011011000"), -- -6.59428e-39 + -7.22511e-39 = -1.38194e-38
	(b"00000000010101000100110010110100", b"00000000000000000000000000000000"),
	(b"00000000010000011100100110011001", b"00000000100101100001011001001101"), -- 7.7417e-39 + 6.04163e-39 = 1.37833e-38
	(b"10000000000010101010111101111110", b"00000000000000000000000000000000"),
	(b"10000000010001010100111100111101", b"10000000010011111111111010111011"), -- -9.8131e-40 + -6.36507e-39 = -7.34638e-39
	(b"00000000011110010100001000100111", b"00000000000000000000000000000000"),
	(b"10000000001111000001110110101001", b"00000000001111010010010001111110"), -- 1.11358e-38 + -5.52077e-39 = 5.61506e-39
	(b"00000000010001111010110001011110", b"00000000000000000000000000000000"),
	(b"10000000000100010110110010100010", b"00000000001101100011111110111100"), -- 6.58215e-39 + -1.60017e-39 = 4.98198e-39
	(b"10000000000100011111101000011011", b"00000000000000000000000000000000"),
	(b"10000000000111111110001110101110", b"10000000001100011101110111001001"), -- -1.65092e-39 + -2.92858e-39 = -4.5795e-39
	(b"10000000010011101110010001101001", b"00000000000000000000000000000000"),
	(b"00000000011000101011011010000010", b"00000000000100111101001000011001"), -- -7.24511e-39 + 9.06535e-39 = 1.82024e-39
	(b"00000000000001111010000101110011", b"00000000000000000000000000000000"),
	(b"00000000001100001011000011100111", b"00000000001110000101001001011010"), -- 7.00766e-40 + 4.47156e-39 = 5.17233e-39
	(b"00000000011001001101111001100101", b"00000000000000000000000000000000"),
	(b"00000000000001100101100001011010", b"00000000011010110011011010111111"), -- 9.26333e-39 + 5.82708e-40 = 9.84604e-39
	(b"10000000000010001110000000100001", b"00000000000000000000000000000000"),
	(b"00000000001110000001001110100000", b"00000000001011110011001101111111"), -- -8.15086e-40 + 5.14983e-39 = 4.33474e-39
	(b"00000000000100110000100100000100", b"00000000000000000000000000000000"),
	(b"00000000000000110111001000111010", b"00000000000101100111101100111110"), -- 1.74811e-39 + 3.16483e-40 = 2.06459e-39
	(b"00000000011100011101101001010110", b"00000000000000000000000000000000"),
	(b"10000000011010101011100011111010", b"00000000000001110010000101011100"), -- 1.04557e-38 + -9.80092e-39 = 6.54816e-40
	(b"10000000001010110101101010000110", b"00000000000000000000000000000000"),
	(b"10000000011001101111011000000110", b"10000000100100100101000010001100"), -- -3.9814e-39 + -9.45548e-39 = -1.34369e-38
	(b"10000000011101010111110110010011", b"00000000000000000000000000000000"),
	(b"10000000011000100001000011000000", b"10000000110101111000111001010011"), -- -1.07898e-38 + -9.00589e-39 = -1.97957e-38
	(b"00000000011000001010000011100000", b"00000000000000000000000000000000"),
	(b"10000000001110111101111110101010", b"00000000001001001100000100110110"), -- 8.87392e-39 + -5.49853e-39 = 3.37539e-39
	(b"00000000011000010110010000110010", b"00000000000000000000000000000000"),
	(b"00000000011011010101011110110010", b"00000000110011101011101111100100"), -- 8.94399e-39 + 1.00415e-38 = 1.89855e-38
	(b"10000000011000000101000111101100", b"00000000000000000000000000000000"),
	(b"10000000010010010100011111100001", b"10000000101010011001100111001101"), -- -8.8456e-39 + -6.72978e-39 = -1.55754e-38
	(b"10000000010110011101010011101110", b"00000000000000000000000000000000"),
	(b"00000000010101011011011101101011", b"10000000000001000001110110000011"), -- -8.24974e-39 + 7.87182e-39 = -3.77929e-40
	(b"00000000011000111100100111001001", b"00000000000000000000000000000000"),
	(b"00000000001110111001011111110111", b"00000000100111110110000111000000"), -- 9.1641e-39 + 5.47281e-39 = 1.46369e-38
	(b"00000000001010010001011001110010", b"00000000000000000000000000000000"),
	(b"00000000000011111110100110010010", b"00000000001110010000000000000100"), -- 3.77331e-39 + 1.46132e-39 = 5.23463e-39
	(b"00000000000010101001100001001010", b"00000000000000000000000000000000"),
	(b"10000000000010111100001101000101", b"10000000000000010010101011111011"), -- 9.72986e-40 + -1.08024e-39 = -1.07254e-40
	(b"10000000011110000011001111001001", b"00000000000000000000000000000000"),
	(b"00000000001100101101100110011100", b"10000000010001010101101000101101"), -- -1.10388e-38 + 4.66984e-39 = -6.369e-39
	(b"10000000000001100101000001111001", b"00000000000000000000000000000000"),
	(b"10000000001000101011111011100110", b"10000000001010010000111101011111"), -- -5.79881e-40 + -3.19089e-39 = -3.77077e-39
	(b"10000000001100010010010010010111", b"00000000000000000000000000000000"),
	(b"10000000001101010101001100111111", b"10000000011001100111011111010110"), -- -4.51307e-39 + -4.89714e-39 = -9.41021e-39
	(b"00000000000001000010100100010100", b"00000000000000000000000000000000"),
	(b"00000000010001010011010000101110", b"00000000010010010101110101000010"), -- 3.82078e-40 + 6.35537e-39 = 6.73745e-39
	(b"00000000010101111110000011110001", b"00000000000000000000000000000000"),
	(b"10000000000111001100110001011001", b"00000000001110110001010010011000"), -- 8.07038e-39 + -2.6447e-39 = 5.42568e-39
	(b"00000000001010110101101110111100", b"00000000000000000000000000000000"),
	(b"00000000001011101010101101101011", b"00000000010110100000011100100111"), -- 3.98183e-39 + 4.28593e-39 = 8.26776e-39
	(b"10000000011111100110111001111111", b"00000000000000000000000000000000"),
	(b"10000000001000111000100101010001", b"10000000101000011111011111010000"), -- -1.16109e-38 + -3.2635e-39 = -1.48744e-38
	(b"00000000010011101100001111111000", b"00000000000000000000000000000000"),
	(b"00000000010010101010110101010111", b"00000000100110010111000101001111"), -- 7.23347e-39 + 6.85801e-39 = 1.40915e-38
	(b"00000000001101110010100001101001", b"00000000000000000000000000000000"),
	(b"10000000000010110000011111101111", b"00000000001011000010000001111010"), -- 5.06545e-39 + -1.01304e-39 = 4.05241e-39
	(b"00000000000000110011011100000111", b"00000000000000000000000000000000"),
	(b"00000000011100101101001101010010", b"00000000011101100000101001011001"), -- 2.95247e-40 + 1.05451e-38 = 1.08403e-38
	(b"00000000011110011111110001111110", b"00000000000000000000000000000000"),
	(b"00000000000110101100110000110100", b"00000000100101001100100010110010"), -- 1.12027e-38 + 2.46098e-39 = 1.36636e-38
	(b"10000000001110011001100110111101", b"00000000000000000000000000000000"),
	(b"10000000010010011111010001110000", b"10000000100000111000111000101101"), -- -5.28977e-39 + -6.79168e-39 = -1.20815e-38
	(b"10000000001011110110011011100110", b"00000000000000000000000000000000"),
	(b"00000000011011111001100011011110", b"00000000010000000011000111111000"), -- -4.35318e-39 + 1.02486e-38 = 5.8954e-39
	(b"10000000001001001011110101110000", b"00000000000000000000000000000000"),
	(b"00000000001111010000110001011010", b"00000000000110000100111011101010"), -- -3.37404e-39 + 5.6064e-39 = 2.23236e-39
	(b"10000000000010111111111110000010", b"00000000000000000000000000000000"),
	(b"00000000010011011101011110110001", b"00000000010000011101100000101111"), -- -1.10185e-39 + 7.14871e-39 = 6.04686e-39
	(b"00000000010010101110001000000101", b"00000000000000000000000000000000"),
	(b"00000000001100011010000010000011", b"00000000011111001000001010001000"), -- 6.87691e-39 + 4.55752e-39 = 1.14344e-38
	(b"10000000010101111000101101010010", b"00000000000000000000000000000000"),
	(b"00000000001101100101000110001010", b"10000000001000010011100111001000"), -- -8.03967e-39 + 4.98837e-39 = -3.0513e-39
	(b"10000000010111010011101110100000", b"00000000000000000000000000000000"),
	(b"00000000010101001101000110100101", b"10000000000010000110100111111011"), -- -8.56209e-39 + 7.78939e-39 = -7.72703e-40
	(b"10000000000011001110101101110100", b"00000000000000000000000000000000"),
	(b"10000000011010111010000101010101", b"10000000011110001000110011001001"), -- -1.18649e-39 + -9.88427e-39 = -1.10708e-38
	(b"10000000001010101010011110011101", b"00000000000000000000000000000000"),
	(b"00000000000000100000000010001101", b"10000000001010001010011100010000"), -- -3.91722e-39 + 1.83869e-40 = -3.73335e-39
	(b"10000000010100001000010100110100", b"00000000000000000000000000000000"),
	(b"00000000011100111001001000010100", b"00000000001000110000110011100000"), -- -7.39462e-39 + 1.06135e-38 = 3.21886e-39
	(b"10000000010100001000010101100010", b"00000000000000000000000000000000"),
	(b"10000000011011101110100100001111", b"10000000101111110110111001110001"), -- -7.39469e-39 + -1.01855e-38 = -1.75802e-38
	(b"10000000011010101100011000010001", b"00000000000000000000000000000000"),
	(b"10000000001111000111001011001011", b"10000000101001110011100011011100"), -- -9.80562e-39 + -5.55131e-39 = -1.53569e-38
	(b"10000000000100000010011001001101", b"00000000000000000000000000000000"),
	(b"10000000010110010010001100000101", b"10000000011010010100100101010010"), -- -1.48311e-39 + -8.18592e-39 = -9.66903e-39
	(b"10000000010111000100000111110010", b"00000000000000000000000000000000"),
	(b"10000000011110101111011111111110", b"10000000110101110011100111110000"), -- -8.47252e-39 + -1.12929e-38 = -1.97654e-38
	(b"10000000010111111011000100000110", b"00000000000000000000000000000000"),
	(b"00000000001011000010101010011011", b"10000000001100111000011001101011"), -- -8.78788e-39 + 4.05605e-39 = -4.73183e-39
	(b"10000000010100111111110111001111", b"00000000000000000000000000000000"),
	(b"10000000001101001001111110000001", b"10000000100010001001110101010000"), -- -7.7134e-39 + -4.83267e-39 = -1.25461e-38
	(b"00000000001000110000101010101010", b"00000000000000000000000000000000"),
	(b"10000000011010000001101011111111", b"10000000010001010001000001010101"), -- 3.21807e-39 + -9.56058e-39 = -6.34251e-39
	(b"10000000010111011010100111111100", b"00000000000000000000000000000000"),
	(b"00000000010110100011100110001011", b"10000000000000110111000001110001"), -- -8.60168e-39 + 8.28584e-39 = -3.15843e-40
	(b"10000000011010100010111001000100", b"00000000000000000000000000000000"),
	(b"10000000001111010111111010101100", b"10000000101001111010110011110000"), -- -9.75116e-39 + -5.64741e-39 = -1.53986e-38
	(b"00000000010110001000001000001000", b"00000000000000000000000000000000"),
	(b"10000000001011001011010100010000", b"00000000001010111100110011111000"), -- 8.12817e-39 + -4.10571e-39 = 4.02246e-39
	(b"10000000000111111101101100110001", b"00000000000000000000000000000000"),
	(b"10000000011000011111011101110100", b"10000000100000011101001010100101"), -- -2.92553e-39 + -8.99681e-39 = -1.19223e-38
	(b"10000000001100000110011010000111", b"00000000000000000000000000000000"),
	(b"00000000010110111101110011011111", b"00000000001010110111011001011000"), -- -4.44488e-39 + 8.43626e-39 = 3.99138e-39
	(b"00000000010010110000100011011010", b"00000000000000000000000000000000"),
	(b"10000000001011111001011100011101", b"00000000000110110111000110111101"), -- 6.89084e-39 + -4.37048e-39 = 2.52036e-39
	(b"10000000011000000010001000000000", b"00000000000000000000000000000000"),
	(b"10000000011001010000111100110010", b"10000000110001010011000100110010"), -- -8.8284e-39 + -9.28084e-39 = -1.81092e-38
	(b"00000000001000000100010101000000", b"00000000000000000000000000000000"),
	(b"10000000010101100000010010000011", b"10000000001101011011111101000011"), -- 2.96358e-39 + -7.89947e-39 = -4.93589e-39
	(b"00000000010011110000110101010000", b"00000000000000000000000000000000"),
	(b"10000000000010111001011100111101", b"00000000010000110111011000010011"), -- 7.25978e-39 + -1.06444e-39 = 6.19534e-39
	(b"10000000011001110000101001000010", b"00000000000000000000000000000000"),
	(b"10000000011001010000100101100101", b"10000000110011000001001110100111"), -- -9.46274e-39 + -9.27876e-39 = -1.87415e-38
	(b"00000000001011100000110101010001", b"00000000000000000000000000000000"),
	(b"10000000011110111011101100011100", b"10000000010011011010110111001011"), -- 4.22921e-39 + -1.13629e-38 = -7.13368e-39
	(b"10000000000000100101011110010101", b"00000000000000000000000000000000"),
	(b"00000000000100100010101100010010", b"00000000000011111101001101111101"), -- -2.1509e-40 + 1.66849e-39 = 1.4534e-39
	(b"00000000001011100101001000000010", b"00000000000000000000000000000000"),
	(b"10000000011001101001100111001000", b"10000000001110000100011111000110"), -- 4.25385e-39 + -9.42239e-39 = -5.16854e-39
	(b"10000000010011100100110001110001", b"00000000000000000000000000000000"),
	(b"10000000000011101000110010001011", b"10000000010111001101100011111100"), -- -7.19059e-39 + -1.33611e-39 = -8.5267e-39
	(b"10000000001110110001111111001011", b"00000000000000000000000000000000"),
	(b"10000000000011011000010010100011", b"10000000010010001010010001101110"), -- -5.4297e-39 + -1.24144e-39 = -6.67114e-39
	(b"10000000000100111011000010000111", b"00000000000000000000000000000000"),
	(b"00000000010101111001011001100000", b"00000000010000111110010111011001"), -- -1.8082e-39 + 8.04363e-39 = 6.23543e-39
	(b"00000000010001011011101101010101", b"00000000000000000000000000000000"),
	(b"00000000001010100101101011000011", b"00000000011100000001011000011000"), -- 6.40385e-39 + 3.88965e-39 = 1.02935e-38
	(b"00000000011101110011101100111110", b"00000000000000000000000000000000"),
	(b"00000000000101111100000101011101", b"00000000100011101111110010011011"), -- 1.09497e-38 + 2.18158e-39 = 1.31313e-38
	(b"00000000000100101011111111010111", b"00000000000000000000000000000000"),
	(b"10000000010011111111011001111100", b"10000000001111010011011010100101"), -- 1.72186e-39 + -7.34343e-39 = -5.62157e-39
	(b"00000000000010111010101001110011", b"00000000000000000000000000000000"),
	(b"00000000011100111001101000001011", b"00000000011111110100010001111110"), -- 1.07134e-39 + 1.06163e-38 = 1.16877e-38
	(b"00000000011011100110001010110010", b"00000000000000000000000000000000"),
	(b"10000000000011011001110010000101", b"00000000011000001100011000101101"), -- 1.01373e-38 + -1.25001e-39 = 8.8873e-39
	(b"10000000001111001100101111000100", b"00000000000000000000000000000000"),
	(b"00000000010011100001111110111010", b"00000000000100010101001111110110"), -- -5.58323e-39 + 7.17455e-39 = 1.59132e-39
	(b"00000000001110000000101001011110", b"00000000000000000000000000000000"),
	(b"10000000001101011001010100011111", b"00000000000000100111010100111111"), -- 5.14651e-39 + -4.92078e-39 = 2.25731e-40
	(b"00000000010100100111011010011000", b"00000000000000000000000000000000"),
	(b"00000000010011101010001111000001", b"00000000101000010001101001011001"), -- 7.57305e-39 + 7.22191e-39 = 1.4795e-38
	(b"10000000001110100111000101111100", b"00000000000000000000000000000000"),
	(b"10000000000000000011101100100110", b"10000000001110101010110010100010"), -- -5.36717e-39 + -2.12185e-41 = -5.38839e-39
	(b"00000000011101101100101100110010", b"00000000000000000000000000000000"),
	(b"10000000011110001110001101100111", b"10000000000000100001100000110101"), -- 1.09095e-38 + -1.11018e-38 = -1.92355e-40
	(b"00000000010111010110001011110100", b"00000000000000000000000000000000"),
	(b"10000000010000010101111110100101", b"00000000000111000000001101001111"), -- 8.5762e-39 + -6.00362e-39 = 2.57258e-39
	(b"00000000000011001110010000010011", b"00000000000000000000000000000000"),
	(b"00000000001001100110110001000111", b"00000000001100110101000001011010"), -- 1.18384e-39 + 3.52859e-39 = 4.71244e-39
	(b"00000000011001101011101111001000", b"00000000000000000000000000000000"),
	(b"10000000000010110111011000011011", b"00000000010110110100010110101101"), -- 9.43458e-39 + -1.05256e-39 = 8.38203e-39
	(b"10000000001010000101101100010010", b"00000000000000000000000000000000"),
	(b"00000000001001110100011110001111", b"10000000000000010001001110000011"), -- -3.70609e-39 + 3.60725e-39 = -9.8835e-41
	(b"00000000010110010000000010000000", b"00000000000000000000000000000000"),
	(b"00000000010001000001010000111100", b"00000000100111010001010010111100"), -- 8.17354e-39 + 6.25207e-39 = 1.44256e-38
	(b"10000000011000000111001011100111", b"00000000000000000000000000000000"),
	(b"10000000010100111000101100111111", b"10000000101100111111111000100110"), -- -8.85743e-39 + -7.6723e-39 = -1.65297e-38
	(b"10000000001010011110001011100100", b"00000000000000000000000000000000"),
	(b"10000000010101010011001101111011", b"10000000011111110001011001011111"), -- -3.84665e-39 + -7.82448e-39 = -1.16711e-38
	(b"00000000011010111100000000011110", b"00000000000000000000000000000000"),
	(b"10000000011011001000100110011000", b"10000000000000001100100101111010"), -- 9.89532e-39 + -9.96759e-39 = -7.22762e-41
	(b"10000000000000001011110001111110", b"00000000000000000000000000000000"),
	(b"00000000010011111000100011001010", b"00000000010011101100110001001100"), -- -6.76183e-41 + 7.30407e-39 = 7.23646e-39
	(b"10000000001101011001010011110110", b"00000000000000000000000000000000"),
	(b"00000000000001000011010010100100", b"10000000001100010110000001010010"), -- -4.92072e-39 + 3.86226e-40 = -4.53449e-39
	(b"00000000001010000011000011010000", b"00000000000000000000000000000000"),
	(b"00000000010010010000011110111110", b"00000000011100010011100010001110"), -- 3.69093e-39 + 6.70677e-39 = 1.03977e-38
	(b"10000000001011010101011010101100", b"00000000000000000000000000000000"),
	(b"10000000011010011110101001101101", b"10000000100101110100000100011001"), -- -4.16369e-39 + -9.72682e-39 = -1.38905e-38
	(b"10000000011000010100100111000110", b"00000000000000000000000000000000"),
	(b"10000000000000010011101100101001", b"10000000011000101000010011101111"), -- -8.93451e-39 + -1.13058e-40 = -9.04757e-39
	(b"00000000010000100010001100001000", b"00000000000000000000000000000000"),
	(b"00000000010010100001101011111110", b"00000000100011000011111000000110"), -- 6.07371e-39 + 6.80551e-39 = 1.28792e-38
	(b"10000000011000000110010011110001", b"00000000000000000000000000000000"),
	(b"10000000010110111011000001010010", b"10000000101111000001010101000011"), -- -8.85242e-39 + -8.42028e-39 = -1.72727e-38
	(b"00000000000000001101110100010100", b"00000000000000000000000000000000"),
	(b"10000000001111110001111110001111", b"10000000001111100100001001111011"), -- 7.93079e-41 + -5.79696e-39 = -5.71765e-39
	(b"10000000010000111010101001001010", b"00000000000000000000000000000000"),
	(b"00000000001110111010100110011100", b"10000000000010000000000010101110"), -- -6.21407e-39 + 5.47914e-39 = -7.34928e-40
	(b"00000000000010100010001010110000", b"00000000000000000000000000000000"),
	(b"10000000010111011000011001111101", b"10000000010100110110001111001101"), -- 9.30798e-40 + -8.58895e-39 = -7.65815e-39
	(b"00000000000100110010100100110011", b"00000000000000000000000000000000"),
	(b"10000000010110001110000001000010", b"10000000010001011011011100001111"), -- 1.75965e-39 + -8.16197e-39 = -6.40232e-39
	(b"00000000010110111010110000010000", b"00000000000000000000000000000000"),
	(b"10000000011011110000000001010100", b"10000000000100110101010001000100"), -- 8.41875e-39 + -1.01939e-38 = -1.7751e-39
	(b"00000000010000011000101011100000", b"00000000000000000000000000000000"),
	(b"10000000010101001100011000110101", b"10000000000100110011101101010101"), -- 6.01913e-39 + -7.78528e-39 = -1.76616e-39
	(b"00000000010110010010011100011101", b"00000000000000000000000000000000"),
	(b"10000000010011011100100100011000", b"00000000000010110101111000000101"), -- 8.18739e-39 + -7.14347e-39 = 1.04392e-39
	(b"10000000000000011101110110111101", b"00000000000000000000000000000000"),
	(b"10000000000001010110111101000001", b"10000000000001110100110011111110"), -- -1.7138e-40 + -4.99088e-40 = -6.70468e-40
	(b"00000000000111001100110100111001", b"00000000000000000000000000000000"),
	(b"00000000011100101111110110001001", b"00000000100011111100101011000010"), -- 2.64501e-39 + 1.05602e-38 = 1.32052e-38
	(b"00000000001010001011010110011100", b"00000000000000000000000000000000"),
	(b"00000000011111011110101010001111", b"00000000101001101010000000101011"), -- 3.73857e-39 + 1.15636e-38 = 1.53021e-38
	(b"10000000011011100010101110011100", b"00000000000000000000000000000000"),
	(b"00000000011000011010110100100100", b"10000000000011000111111001111000"), -- -1.01175e-38 + 8.97015e-39 = -1.14739e-39
	(b"00000000000001111100000101000011", b"00000000000000000000000000000000"),
	(b"00000000010111110101010110100110", b"00000000011001110001011011101001"), -- 7.12178e-40 + 8.7551e-39 = 9.46727e-39
	(b"00000000011010011101100110001000", b"00000000000000000000000000000000"),
	(b"10000000000110011101100111011001", b"00000000010011111111111110101111"), -- 9.72076e-39 + -2.37404e-39 = 7.34673e-39
	(b"00000000010101001001001010010101", b"00000000000000000000000000000000"),
	(b"00000000011010011001100100011101", b"00000000101111100010101110110010"), -- 7.76677e-39 + 9.69765e-39 = 1.74644e-38
	(b"00000000001101010011110001100011", b"00000000000000000000000000000000"),
	(b"00000000011101010100010011100110", b"00000000101010101000000101001001"), -- 4.88894e-39 + 1.07695e-38 = 1.56584e-38
	(b"00000000001101100011110100110110", b"00000000000000000000000000000000"),
	(b"10000000000101100100110010010110", b"00000000000111111111000010100000"), -- 4.98108e-39 + -2.04785e-39 = 2.93322e-39
	(b"00000000001001111111011001011110", b"00000000000000000000000000000000"),
	(b"00000000000111000000101000010010", b"00000000010001000000000001110000"), -- 3.66996e-39 + 2.57501e-39 = 6.24497e-39
	(b"10000000001001010101010101101010", b"00000000000000000000000000000000"),
	(b"10000000000101101110101010110111", b"10000000001111000100000000100001"), -- -3.42855e-39 + -2.10458e-39 = -5.53313e-39
	(b"00000000011001110110101100010000", b"00000000000000000000000000000000"),
	(b"00000000000110111011011100100000", b"00000000100000110010001000110000"), -- 9.49746e-39 + 2.54525e-39 = 1.20427e-38
	(b"00000000011111100001111001001101", b"00000000000000000000000000000000"),
	(b"10000000011100010100011101111110", b"00000000000011001101011011001111"), -- 1.15821e-38 + -1.04031e-38 = 1.17908e-39
	(b"00000000011011010111001000000010", b"00000000000000000000000000000000"),
	(b"10000000001011100110010100011001", b"00000000001111110000110011101001"), -- 1.0051e-38 + -4.2607e-39 = 5.79027e-39
	(b"00000000001001111010101110010111", b"00000000000000000000000000000000"),
	(b"00000000011000101100101111100111", b"00000000100010100111011101111110"), -- 3.64314e-39 + 9.07303e-39 = 1.27162e-38
	(b"00000000001001000111111010011000", b"00000000000000000000000000000000"),
	(b"10000000000000100011010001011100", b"00000000001000100100101000111100"), -- 3.35149e-39 + -2.02454e-40 = 3.14904e-39
	(b"00000000001100010011100011101110", b"00000000000000000000000000000000"),
	(b"00000000000111110010001011010000", b"00000000010100000101101110111110"), -- 4.52036e-39 + 2.85939e-39 = 7.37975e-39
	(b"10000000000111010010000110011000", b"00000000000000000000000000000000"),
	(b"10000000010111010111001100010001", b"10000000011110101001010010101001"), -- -2.67528e-39 + -8.58198e-39 = -1.12573e-38
	(b"00000000001010111001101100000010", b"00000000000000000000000000000000"),
	(b"10000000011100010000011111110001", b"10000000010001010110110011101111"), -- 4.00453e-39 + -1.03803e-38 = -6.37573e-39
	(b"10000000000011001011101111011110", b"00000000000000000000000000000000"),
	(b"10000000001011101010000110000110", b"10000000001110110101110101100100"), -- -1.16942e-39 + -4.28238e-39 = -5.4518e-39
	(b"00000000000100011011011001101001", b"00000000000000000000000000000000"),
	(b"10000000010101101111111000011111", b"10000000010001010100011110110110"), -- 1.62664e-39 + -7.98901e-39 = -6.36237e-39
	(b"10000000011011010001001001100011", b"00000000000000000000000000000000"),
	(b"00000000011001111011000010010100", b"10000000000001010110000111001111"), -- -1.00167e-38 + 9.5224e-39 = -4.94265e-40
	(b"10000000001110000011011011001010", b"00000000000000000000000000000000"),
	(b"00000000001101111011011010011111", b"10000000000000001000000000101011"), -- -5.16244e-39 + 5.11646e-39 = -4.5978e-41
	(b"00000000000111101011000011000000", b"00000000000000000000000000000000"),
	(b"00000000000110011101011000110110", b"00000000001110001000011011110110"), -- 2.81847e-39 + 2.37273e-39 = 5.1912e-39
	(b"10000000010000011001111101011100", b"00000000000000000000000000000000"),
	(b"00000000011110111111110101101011", b"00000000001110100101111000001111"), -- -6.02647e-39 + 1.13867e-38 = 5.3602e-39
	(b"00000000000111001100000010110101", b"00000000000000000000000000000000"),
	(b"00000000000010110110101110111001", b"00000000001010000010110001101110"), -- 2.64052e-39 + 1.04883e-39 = 3.68936e-39
	(b"10000000011110000011100100110100", b"00000000000000000000000000000000"),
	(b"10000000011001000010101101001101", b"10000000110111000110010010000001"), -- -1.10408e-38 + -9.19908e-39 = -2.02399e-38
	(b"00000000011010100001101111101010", b"00000000000000000000000000000000"),
	(b"10000000000011101101011100110100", b"00000000010110110100010010110110"), -- 9.74458e-39 + -1.3629e-39 = 8.38168e-39
	(b"00000000001001011010011011000111", b"00000000000000000000000000000000"),
	(b"10000000000110100111010100111010", b"00000000000010110011000110001101"), -- 3.45774e-39 + -2.42978e-39 = 1.02797e-39
	(b"10000000011011000101000000001100", b"00000000000000000000000000000000"),
	(b"00000000001000110010101010001000", b"10000000010010010010010110000100"), -- -9.94695e-39 + 3.2295e-39 = -6.71745e-39
	(b"00000000010011010011001101101001", b"00000000000000000000000000000000"),
	(b"10000000000001000101110110010010", b"00000000010010001101010111010111"), -- 7.08978e-39 + -4.00909e-40 = 6.68887e-39
	(b"10000000011100001001011001111010", b"00000000000000000000000000000000"),
	(b"00000000000111110110001010101110", b"10000000010100010011001111001100"), -- -1.03396e-38 + 2.8823e-39 = -7.45726e-39
	(b"00000000010101000011011011010001", b"00000000000000000000000000000000"),
	(b"10000000011101010110011100011111", b"10000000001000010011000001001110"), -- 7.73385e-39 + -1.07817e-38 = -3.0479e-39
	(b"00000000000110011000011010000101", b"00000000000000000000000000000000"),
	(b"00000000011010001110111100111101", b"00000000100000100111010111000010"), -- 2.34414e-39 + 9.63671e-39 = 1.19809e-38
	(b"10000000001011000110010001000111", b"00000000000000000000000000000000"),
	(b"00000000000010001010011001100100", b"10000000001000111011110111100011"), -- -4.07673e-39 + 7.94374e-40 = -3.28236e-39
	(b"10000000001101001010011100001000", b"00000000000000000000000000000000"),
	(b"00000000001100110100010101111010", b"10000000000000010110000110001110"), -- -4.83537e-39 + 4.70853e-39 = -1.26832e-40
	(b"10000000000111111001010010110010", b"00000000000000000000000000000000"),
	(b"00000000000100011110100011001101", b"10000000000011011010101111100101"), -- -2.90024e-39 + 1.64472e-39 = -1.25553e-39
	(b"10000000010001111001101101000110", b"00000000000000000000000000000000"),
	(b"10000000011001110011001110100011", b"10000000101011101100111011101001"), -- -6.57602e-39 + -9.47758e-39 = -1.60536e-38
	(b"00000000010010110000101101011100", b"00000000000000000000000000000000"),
	(b"10000000001101101111111100101100", b"00000000000101000000110000110000"), -- 6.89174e-39 + -5.05066e-39 = 1.84108e-39
	(b"10000000000011111100101111001101", b"00000000000000000000000000000000"),
	(b"10000000011001011100000101101101", b"10000000011101011000110100111010"), -- -1.45064e-39 + -9.34477e-39 = -1.07954e-38
	(b"00000000010000001011110100000001", b"00000000000000000000000000000000"),
	(b"00000000010001001011011111111111", b"00000000100001010111010100000000"), -- 5.94527e-39 + 6.31082e-39 = 1.22561e-38
	(b"10000000010111110001101011000011", b"00000000000000000000000000000000"),
	(b"10000000000101011001010011111011", b"10000000011101001010111110111110"), -- -8.73397e-39 + -1.98199e-39 = -1.0716e-38
	(b"10000000001010100100101000011111", b"00000000000000000000000000000000"),
	(b"00000000010000101001001010110011", b"00000000000110000100100010010100"), -- -3.88368e-39 + 6.11377e-39 = 2.23009e-39
	(b"10000000010001111011100010100111", b"00000000000000000000000000000000"),
	(b"10000000001001001010110011111011", b"10000000011011000110010110100010"), -- -6.58656e-39 + -3.36813e-39 = -9.95469e-39
	(b"10000000011100001011111111010001", b"00000000000000000000000000000000"),
	(b"10000000001100011110011100111001", b"10000000101000101010011100001010"), -- -1.03544e-38 + -4.58289e-39 = -1.49373e-38
	(b"10000000011011101010110111101011", b"00000000000000000000000000000000"),
	(b"00000000010101111010001000001011", b"10000000000101110000101111100000"), -- -1.01643e-38 + 8.04782e-39 = -2.11648e-39
	(b"10000000001100110001010010101010", b"00000000000000000000000000000000"),
	(b"00000000001101001000100010100011", b"00000000000000010111001111111001"), -- -4.69102e-39 + 4.82446e-39 = 1.33439e-40
	(b"00000000001100000100101011110101", b"00000000000000000000000000000000"),
	(b"00000000011011000010101101010110", b"00000000100111000111011001001011"), -- 4.43499e-39 + 9.93378e-39 = 1.43688e-38
	(b"10000000000100101010010000000110", b"00000000000000000000000000000000"),
	(b"10000000001010000011101101010110", b"10000000001110101101111101011100"), -- -1.71188e-39 + -3.69471e-39 = -5.40659e-39
	(b"00000000010111110110110001101100", b"00000000000000000000000000000000"),
	(b"00000000010010011010101110100000", b"00000000101010010001100000001100"), -- 8.76327e-39 + 6.76556e-39 = 1.55288e-38
	(b"10000000000001101101101111001001", b"00000000000000000000000000000000"),
	(b"10000000011111011010011000001111", b"10000000100001001000000111011000"), -- -6.29857e-40 + -1.1539e-38 = -1.21689e-38
	(b"00000000001011000000010011011011", b"00000000000000000000000000000000"),
	(b"00000000010101011110110001000010", b"00000000100000011111000100011101"), -- 4.0425e-39 + 7.89077e-39 = 1.19333e-38
	(b"10000000010000001100001000010010", b"00000000000000000000000000000000"),
	(b"10000000000010110101001111100010", b"10000000010011000001010111110100"), -- -5.94709e-39 + -1.04028e-39 = -6.98737e-39
	(b"00000000011101110011001111010011", b"00000000000000000000000000000000"),
	(b"00000000010010101011011001101001", b"00000000110000011110101000111100"), -- 1.0947e-38 + 6.86126e-39 = 1.78083e-38
	(b"00000000001110010101100011001000", b"00000000000000000000000000000000"),
	(b"10000000011100000100010100110011", b"10000000001101101110110001101011"), -- 5.26647e-39 + -1.03104e-38 = -5.04393e-39
	(b"10000000001100101000010110010001", b"00000000000000000000000000000000"),
	(b"10000000010110000000001111010100", b"10000000100010101000100101100101"), -- -4.63969e-39 + -8.0829e-39 = -1.27226e-38
	(b"10000000001101001100100000101110", b"00000000000000000000000000000000"),
	(b"10000000011100100110111100010001", b"10000000101001110011011100111111"), -- -4.84726e-39 + -1.05091e-38 = -1.53563e-38
	(b"00000000011101000100001010001010", b"00000000000000000000000000000000"),
	(b"10000000010010010011110000101111", b"00000000001010110000011001011011"), -- 1.06768e-38 + -6.72558e-39 = 3.95121e-39
	(b"10000000001101111010001111111101", b"00000000000000000000000000000000"),
	(b"00000000010100111101010000010010", b"00000000000111000011000000010101"), -- -5.10978e-39 + 7.69842e-39 = 2.58864e-39
	(b"10000000010001101010100101011010", b"00000000000000000000000000000000"),
	(b"00000000000001000000110011001111", b"10000000010000101001110010001011"), -- -6.48924e-39 + 3.71937e-40 = -6.1173e-39
	(b"10000000010111001111110101101110", b"00000000000000000000000000000000"),
	(b"00000000011111001011011001100001", b"00000000000111111011100011110011"), -- -8.53978e-39 + 1.1453e-38 = 2.91325e-39
	(b"10000000000001111110110101010111", b"00000000000000000000000000000000"),
	(b"00000000000101110001100000110110", b"00000000000011110010101011011111"), -- -7.2799e-40 + 2.1209e-39 = 1.39291e-39
	(b"00000000010001101100010110011000", b"00000000000000000000000000000000"),
	(b"00000000011101110011000010111111", b"00000000101111011111011001010111"), -- 6.49937e-39 + 1.09459e-38 = 1.74453e-38
	(b"10000000001101101000011101010111", b"00000000000000000000000000000000"),
	(b"10000000001010110110011000100000", b"10000000011000011110110101110111"), -- -5.00767e-39 + -3.98556e-39 = -8.99323e-39
	(b"10000000001001100001110010010000", b"00000000000000000000000000000000"),
	(b"00000000001101001110000101110000", b"00000000000011101100010011100000"), -- -3.5e-39 + 4.85632e-39 = 1.35632e-39
	(b"10000000010111111011000110001011", b"00000000000000000000000000000000"),
	(b"00000000001111101101100010001111", b"10000000001000001101100011111100"), -- -8.78806e-39 + 5.77149e-39 = -3.01658e-39
	(b"10000000000000010001010001011111", b"00000000000000000000000000000000"),
	(b"00000000011110100001100100111010", b"00000000011110010000010011011011"), -- -9.91433e-41 + 1.1213e-38 = 1.11138e-38
	(b"10000000011000000101001101101011", b"00000000000000000000000000000000"),
	(b"00000000000010101110110110100110", b"10000000010101010110010111000101"), -- -8.84613e-39 + 1.00361e-39 = -7.84253e-39
	(b"00000000010011100111010011110110", b"00000000000000000000000000000000"),
	(b"00000000010001110001010110001101", b"00000000100101011000101010000011"), -- 7.20513e-39 + 6.52805e-39 = 1.37332e-38
	(b"10000000001110101111101011011101", b"00000000000000000000000000000000"),
	(b"10000000010100000010110111000000", b"10000000100010110010100010011101"), -- -5.41645e-39 + -7.36325e-39 = -1.27797e-38
	(b"00000000000000000100100001100011", b"00000000000000000000000000000000"),
	(b"10000000001111111110110111010101", b"10000000001111111010010101110010"), -- 2.59675e-41 + -5.87095e-39 = -5.84499e-39
	(b"00000000001000011101010100011101", b"00000000000000000000000000000000"),
	(b"10000000001110101011001010010101", b"10000000000110001101110101111000"), -- 3.10702e-39 + -5.39052e-39 = -2.2835e-39
	(b"10000000010101001001100111101000", b"00000000000000000000000000000000"),
	(b"10000000010101111011101011011100", b"10000000101011000101010011000100"), -- -7.76939e-39 + -8.05672e-39 = -1.58261e-38
	(b"10000000000001101100111010101010", b"00000000000000000000000000000000"),
	(b"10000000001010100011011000101011", b"10000000001100010000010011010101"), -- -6.2515e-40 + -3.87652e-39 = -4.50167e-39
	(b"00000000011111100111111111010011", b"00000000000000000000000000000000"),
	(b"00000000001100100000110011011100", b"00000000101100001000110010101111"), -- 1.16171e-38 + 4.59639e-39 = 1.62135e-38
	(b"00000000010100000000010100111000", b"00000000000000000000000000000000"),
	(b"00000000001001010011001011110100", b"00000000011101010011100000101100"), -- 7.34871e-39 + 3.41619e-39 = 1.07649e-38
	(b"10000000000000110100110100110011", b"00000000000000000000000000000000"),
	(b"10000000001101101110101100111011", b"10000000001110100011100001101110"), -- -3.032e-40 + -5.0435e-39 = -5.3467e-39
	(b"10000000010110001101010001111000", b"00000000000000000000000000000000"),
	(b"00000000001010100010110011101010", b"10000000001011101010011110001110"), -- -8.15774e-39 + 3.8732e-39 = -4.28454e-39
	(b"00000000010000010001001010001111", b"00000000000000000000000000000000"),
	(b"10000000000010011110010101011011", b"00000000001101110010110100110100"), -- 5.97596e-39 + -9.08797e-40 = 5.06717e-39
	(b"10000000010010010110101101101010", b"00000000000000000000000000000000"),
	(b"00000000010000001101010111100101", b"10000000000010001001010110000101"), -- -6.74252e-39 + 5.9542e-39 = -7.88321e-40
	(b"00000000011111101100111010001111", b"00000000000000000000000000000000"),
	(b"00000000001001010011000110111001", b"00000000101001000000000001001000"), -- 1.16454e-38 + 3.41575e-39 = 1.50611e-38
	(b"10000000010111100000110101100000", b"00000000000000000000000000000000"),
	(b"00000000000100100111111101011101", b"10000000010010111000111000000011"), -- -8.63733e-39 + 1.69873e-39 = -6.93861e-39
	(b"10000000000010000101010010101101", b"00000000000000000000000000000000"),
	(b"10000000000110000011110000011000", b"10000000001000001001000011000101"), -- -7.6506e-40 + -2.22561e-39 = -2.99067e-39
	(b"10000000001000000111101100001110", b"00000000000000000000000000000000"),
	(b"10000000010011001110101101110011", b"10000000011011010110011010000001"), -- -2.98288e-39 + -7.06396e-39 = -1.00468e-38
	(b"00000000000000010000111100011101", b"00000000000000000000000000000000"),
	(b"00000000011010010010100001100100", b"00000000011010100011011110000001"), -- 9.72571e-41 + 9.65722e-39 = 9.75447e-39
	(b"10000000001101001000001101010101", b"00000000000000000000000000000000"),
	(b"00000000010100000001001101001000", b"00000000000110111000111111110011"), -- -4.82256e-39 + 7.35376e-39 = 2.5312e-39
	(b"00000000011000011010000100011110", b"00000000000000000000000000000000"),
	(b"10000000000100000101000111111000", b"00000000010100010100111100100110"), -- 8.96584e-39 + -1.49877e-39 = 7.46707e-39
	(b"10000000010110011000011001001111", b"00000000000000000000000000000000"),
	(b"10000000000110010101111010000000", b"10000000011100101110010011001111"), -- -8.22154e-39 + -2.32979e-39 = -1.05513e-38
	(b"10000000001101101100000010010011", b"00000000000000000000000000000000"),
	(b"10000000010110000110110101101000", b"10000000100011110010110111111011"), -- -5.0282e-39 + -8.12077e-39 = -1.3149e-38
	(b"10000000000010100111111100001110", b"00000000000000000000000000000000"),
	(b"10000000000111010110000111001101", b"10000000001001111110000011011011"), -- -9.63934e-40 + -2.69831e-39 = -3.66225e-39
	(b"00000000001101110000110100111011", b"00000000000000000000000000000000"),
	(b"10000000011100000111110110010110", b"10000000001110010111000001011011"), -- 5.0557e-39 + -1.03306e-38 = -5.27493e-39
	(b"00000000000101010111111110011100", b"00000000000000000000000000000000"),
	(b"00000000010010110010010111011001", b"00000000011000001010010101110101"), -- 1.97432e-39 + 6.90124e-39 = 8.87556e-39
	(b"10000000000010101110110100111100", b"00000000000000000000000000000000"),
	(b"10000000000001111001010111011001", b"10000000000100101000001100010101"), -- -1.00346e-39 + -6.96604e-40 = -1.70006e-39
	(b"00000000001110101110111010010001", b"00000000000000000000000000000000"),
	(b"00000000011101101100011010001000", b"00000000101100011011010100011001"), -- 5.41204e-39 + 1.09078e-38 = 1.63198e-38
	(b"00000000000011010011010101111000", b"00000000000000000000000000000000"),
	(b"00000000000000110110001110010100", b"00000000000100001001100100001100"), -- 1.21304e-39 + 3.11228e-40 = 1.52427e-39
	(b"00000000000110001001110100000111", b"00000000000000000000000000000000"),
	(b"00000000001100110001010111000001", b"00000000010010111011001011001000"), -- 2.26038e-39 + 4.69141e-39 = 6.9518e-39
	(b"10000000011001011001100110010111", b"00000000000000000000000000000000"),
	(b"00000000011001001010110011000011", b"10000000000000001110110011010100"), -- -9.33048e-39 + 9.24552e-39 = -8.49579e-41
	(b"00000000010110110011110111001101", b"00000000000000000000000000000000"),
	(b"00000000010100110010001011011011", b"00000000101011100110000010101000"), -- 8.3792e-39 + 7.63485e-39 = 1.60141e-38
	(b"00000000001000000110110111011000", b"00000000000000000000000000000000"),
	(b"00000000011110101000101100000010", b"00000000100110101111100011011010"), -- 2.97814e-39 + 1.12538e-38 = 1.42319e-38
	(b"10000000010010011101100011111101", b"00000000000000000000000000000000"),
	(b"10000000000111001110000001011011", b"10000000011001101011100101011000"), -- -6.78183e-39 + -2.65188e-39 = -9.43371e-39
	(b"00000000001011001010010000000001", b"00000000000000000000000000000000"),
	(b"10000000001000001000110000111111", b"00000000000011000001011111000010"), -- 4.0996e-39 + -2.98905e-39 = 1.11055e-39
	(b"10000000001011000110010111011011", b"00000000000000000000000000000000"),
	(b"00000000010011000011110001011010", b"00000000000111111101011001111111"), -- -4.0773e-39 + 7.00115e-39 = 2.92385e-39
	(b"00000000011100000101001100001111", b"00000000000000000000000000000000"),
	(b"00000000011110000000000000010110", b"00000000111010000101001100100101"), -- 1.03154e-38 + 1.10203e-38 = 2.13357e-38
	(b"00000000011001000101100101101110", b"00000000000000000000000000000000"),
	(b"10000000011001100110100110011011", b"10000000000000100001000000101101"), -- 9.21563e-39 + -9.4051e-39 = -1.89474e-40
	(b"10000000011001100111011001110001", b"00000000000000000000000000000000"),
	(b"00000000000000111110000001011110", b"10000000011000101001011000010011"), -- -9.40971e-39 + 3.55994e-40 = -9.05372e-39
	(b"10000000011110000110000110101110", b"00000000000000000000000000000000"),
	(b"00000000010010000110011110000111", b"10000000001011111111101000100111"), -- -1.10553e-38 + 6.64929e-39 = -4.40601e-39
	(b"10000000010110001011100011111110", b"00000000000000000000000000000000"),
	(b"10000000010101011111001100000110", b"10000000101011101010110000000100"), -- -8.14789e-39 + -7.8932e-39 = -1.60411e-38
	(b"00000000011001101110111000001011", b"00000000000000000000000000000000"),
	(b"00000000001101110110000011110000", b"00000000100111100100111011111011"), -- 9.45261e-39 + 5.08573e-39 = 1.45383e-38
	(b"00000000000101100110001111101100", b"00000000000000000000000000000000"),
	(b"00000000001011000101010101100100", b"00000000010000101011100101010000"), -- 2.05623e-39 + 4.07139e-39 = 6.12762e-39
	(b"00000000010110100011011000101111", b"00000000000000000000000000000000"),
	(b"10000000001001111001111111010001", b"00000000001100101001011001011110"), -- 8.28463e-39 + -3.63892e-39 = 4.64572e-39
	(b"00000000001101000000111100000101", b"00000000000000000000000000000000"),
	(b"10000000000111111011100110111101", b"00000000000101000101010101001000"), -- 4.78083e-39 + -2.91353e-39 = 1.8673e-39
	(b"00000000010110101010001000101011", b"00000000000000000000000000000000"),
	(b"00000000010111100110101000010011", b"00000000101110010000110000111110"), -- 8.32337e-39 + 8.67059e-39 = 1.6994e-38
	(b"10000000010101001011011001000000", b"00000000000000000000000000000000"),
	(b"10000000011011001000100011001010", b"10000000110000010011111100001010"), -- -7.77956e-39 + -9.9673e-39 = -1.77469e-38
	(b"10000000011000001100100010010010", b"00000000000000000000000000000000"),
	(b"10000000010100110010011111111110", b"10000000101100111111000010010000"), -- -8.88816e-39 + -7.63669e-39 = -1.65249e-38
	(b"10000000011110111111111000010101", b"00000000000000000000000000000000"),
	(b"10000000000111100101110011110010", b"10000000100110100101101100000111"), -- -1.13869e-38 + -2.78841e-39 = -1.41753e-38
	(b"10000000000000100011010010111101", b"00000000000000000000000000000000"),
	(b"10000000010001101011110001101100", b"10000000010010001111000100101001"), -- -2.0259e-40 + -6.49608e-39 = -6.69867e-39
	(b"10000000011111110100100000010110", b"00000000000000000000000000000000"),
	(b"00000000001100100100110011000001", b"10000000010011001111101101010101"), -- -1.1689e-38 + 4.61931e-39 = -7.06966e-39
	(b"10000000001100010000011000110101", b"00000000000000000000000000000000"),
	(b"00000000001110010000100010110110", b"00000000000010000000001010000001"), -- -4.50217e-39 + 5.23775e-39 = 7.35582e-40
	(b"00000000001010010011101000101000", b"00000000000000000000000000000000"),
	(b"00000000000100100011111010101111", b"00000000001110110111100011010111"), -- 3.78612e-39 + 1.67553e-39 = 5.46164e-39
	(b"10000000010101101010000000011111", b"00000000000000000000000000000000"),
	(b"10000000001100111011011111101011", b"10000000100010100101100000001010"), -- -7.95529e-39 + -4.74959e-39 = -1.27049e-38
	(b"00000000001001100110101110100111", b"00000000000000000000000000000000"),
	(b"10000000010010010110000010001100", b"10000000001000101111010011100101"), -- 3.52837e-39 + -6.73863e-39 = -3.21026e-39
	(b"00000000000101010011111011111101", b"00000000000000000000000000000000"),
	(b"10000000001010001110110000010011", b"10000000000100111010110100010110"), -- 1.95114e-39 + -3.75811e-39 = -1.80697e-39
	(b"00000000000000010101101010010001", b"00000000000000000000000000000000"),
	(b"00000000010110010111011001100111", b"00000000010110101101000011111000"), -- 1.24325e-40 + 8.21583e-39 = 8.34016e-39
	(b"00000000010111010001101100110101", b"00000000000000000000000000000000"),
	(b"10000000000101010111001100111011", b"00000000010001111010011111111010"), -- 8.55046e-39 + -1.96988e-39 = 6.58058e-39
	(b"00000000010110101010100001001011", b"00000000000000000000000000000000"),
	(b"00000000000110111000010110001000", b"00000000011101100010110111010011"), -- 8.32557e-39 + 2.52746e-39 = 1.0853e-38
	(b"10000000010101100001110010100001", b"00000000000000000000000000000000"),
	(b"00000000000000101001101010000001", b"10000000010100111000001000100000"), -- -7.90812e-39 + 2.39097e-40 = -7.66903e-39
	(b"00000000010001011000010010100001", b"00000000000000000000000000000000"),
	(b"00000000000010010000110000101001", b"00000000010011101001000011001010"), -- 6.38423e-39 + 8.30882e-40 = 7.21511e-39
	(b"10000000000111000010011101100011", b"00000000000000000000000000000000"),
	(b"00000000010100101000010000100011", b"00000000001101100101110011000000"), -- -2.58552e-39 + 7.57791e-39 = 4.99239e-39
	(b"10000000001111010110100111100110", b"00000000000000000000000000000000"),
	(b"00000000010000111011011001001010", b"00000000000001100100110001100100"), -- -5.63995e-39 + 6.21837e-39 = 5.78417e-40
	(b"10000000011011100010110010001110", b"00000000000000000000000000000000"),
	(b"10000000010010111110001011111101", b"10000000101110100000111110001011"), -- -1.01179e-38 + -6.96909e-39 = -1.7087e-38
	(b"00000000010010110011110111100010", b"00000000000000000000000000000000"),
	(b"00000000011110100101010110001001", b"00000000110001011001001101101011"), -- 6.90986e-39 + 1.12346e-38 = 1.81445e-38
	(b"10000000011111001111010101001100", b"00000000000000000000000000000000"),
	(b"00000000011111000101011001110000", b"10000000000000001001111011011100"), -- -1.14756e-38 + 1.14186e-38 = -5.6988e-41
	(b"10000000011010000100011001110100", b"00000000000000000000000000000000"),
	(b"10000000000100011100101001000110", b"10000000011110100001000010111010"), -- -9.57617e-39 + -1.63377e-39 = -1.12099e-38
	(b"10000000011101110101000111101010", b"00000000000000000000000000000000"),
	(b"00000000001110110010111100010001", b"10000000001111000010001011011001"), -- -1.09578e-38 + 5.43518e-39 = -5.52263e-39
	(b"00000000000001010101000010111011", b"00000000000000000000000000000000"),
	(b"00000000011000110110011101111011", b"00000000011010001011100000110110"), -- 4.88138e-40 + 9.12884e-39 = 9.61697e-39
	(b"00000000000000110111001111110011", b"00000000000000000000000000000000"),
	(b"00000000001000001110101001101101", b"00000000001001000101111001100000"), -- 3.17101e-40 + 3.02283e-39 = 3.33993e-39
	(b"00000000001000000010001000010101", b"00000000000000000000000000000000"),
	(b"10000000001011011000110110111100", b"10000000000011010110101110100111"), -- 2.95096e-39 + -4.18344e-39 = -1.23248e-39
	(b"00000000010000110010000010101001", b"00000000000000000000000000000000"),
	(b"10000000000011111011011011111110", b"00000000001100110110100110101011"), -- 6.16469e-39 + -1.44318e-39 = 4.72152e-39
	(b"00000000000010001110111100100101", b"00000000000000000000000000000000"),
	(b"10000000000011001110101011011111", b"10000000000000111111101110111010"), -- 8.20473e-40 + -1.18628e-39 = -3.65809e-40
	(b"00000000001010011001000100111101", b"00000000000000000000000000000000"),
	(b"00000000011000101001011000100010", b"00000000100011000010011101011111"), -- 3.81736e-39 + 9.05374e-39 = 1.28711e-38
	(b"10000000000001111101001100001111", b"00000000000000000000000000000000"),
	(b"00000000001001010101101101110011", b"00000000000111011000100001100100"), -- -7.18562e-40 + 3.43072e-39 = 2.71216e-39
	(b"10000000001010110010011101010101", b"00000000000000000000000000000000"),
	(b"10000000001011011101010000101010", b"10000000010110001111101101111111"), -- -3.96304e-39 + -4.20871e-39 = -8.17174e-39
	(b"10000000010000110101110101001000", b"00000000000000000000000000000000"),
	(b"00000000011110011000010001111000", b"00000000001101100010011100110000"), -- -6.18644e-39 + 1.11596e-38 = 4.97317e-39
	(b"00000000011100110110100001000110", b"00000000000000000000000000000000"),
	(b"00000000010110000001001001101100", b"00000000110010110111101010110010"), -- 1.05985e-38 + 8.08813e-39 = 1.86866e-38
	(b"00000000001000011001100111100010", b"00000000000000000000000000000000"),
	(b"10000000001101001101100001000110", b"10000000000100110011111001100100"), -- 3.08577e-39 + -4.85303e-39 = -1.76726e-39
	(b"00000000001011110010011111100110", b"00000000000000000000000000000000"),
	(b"00000000000010010101101111110010", b"00000000001110001000001111011000"), -- 4.33058e-39 + 8.59503e-40 = 5.19008e-39
	(b"00000000011101110101101100011001", b"00000000000000000000000000000000"),
	(b"10000000000011100100001100100011", b"00000000011010010001011111110110"), -- 1.09611e-38 + -1.30978e-39 = 9.65132e-39
	(b"00000000010010001001000001101110", b"00000000000000000000000000000000"),
	(b"00000000000000001011100101101110", b"00000000010010010100100111011100"), -- 6.66397e-39 + 6.65196e-41 = 6.73049e-39
	(b"10000000000101011010001000000010", b"00000000000000000000000000000000"),
	(b"00000000001100111000100011011110", b"00000000000111011110011011011100"), -- -1.98666e-39 + 4.73271e-39 = 2.74605e-39
	(b"10000000001100100010111101110110", b"00000000000000000000000000000000"),
	(b"10000000011010100111101001101101", b"10000000100111001010100111100011"), -- -4.6088e-39 + -9.77848e-39 = -1.43873e-38
	(b"00000000011111010101010111101100", b"00000000000000000000000000000000"),
	(b"00000000001010011010110111001001", b"00000000101001110000001110110101"), -- 1.15103e-38 + 3.8276e-39 = 1.53379e-38
	(b"10000000001010001001101010100111", b"00000000000000000000000000000000"),
	(b"10000000011101010110100001010100", b"10000000100111100000001011111011"), -- -3.7289e-39 + -1.07822e-38 = -1.45111e-38
	(b"10000000000000101101110111100011", b"00000000000000000000000000000000"),
	(b"10000000000110110011010110001001", b"10000000000111100001001101101100"), -- -2.63269e-40 + -2.49876e-39 = -2.76203e-39
	(b"00000000001011010110011010001001", b"00000000000000000000000000000000"),
	(b"00000000001110011011101101111101", b"00000000011001110010001000000110"), -- 4.16938e-39 + 5.30188e-39 = 9.47126e-39
	(b"10000000000000101101100010110001", b"00000000000000000000000000000000"),
	(b"00000000001100110011001000101110", b"00000000001100000101100101111101"), -- -2.61405e-40 + 4.70161e-39 = 4.44021e-39
	(b"10000000001010001100110011010011", b"00000000000000000000000000000000"),
	(b"10000000010000000010101100011001", b"10000000011010001111011111101100"), -- -3.7469e-39 + -5.89293e-39 = -9.63983e-39
	(b"10000000010110001010111011111110", b"00000000000000000000000000000000"),
	(b"00000000000010101011111000001010", b"10000000010011011111000011110100"), -- -8.1443e-39 + 9.86528e-40 = -7.15777e-39
	(b"00000000011010100001110000010111", b"00000000000000000000000000000000"),
	(b"00000000001111001000010101110111", b"00000000101001101010000110001110"), -- 9.74464e-39 + 5.55801e-39 = 1.53026e-38
	(b"10000000001100110010010000010101", b"00000000000000000000000000000000"),
	(b"10000000001010011100111001000000", b"10000000010111001111001001010101"), -- -4.69655e-39 + -3.83924e-39 = -8.5358e-39
	(b"00000000000111001110000110101101", b"00000000000000000000000000000000"),
	(b"00000000001011001000000100111011", b"00000000010010010110001011101000"), -- 2.65235e-39 + 4.08712e-39 = 6.73947e-39
	(b"00000000001011110000011100011000", b"00000000000000000000000000000000"),
	(b"00000000011011111001101111000001", b"00000000100111101010001011011001"), -- 4.31881e-39 + 1.02496e-38 = 1.45684e-38
	(b"00000000001010111101101011111111", b"00000000000000000000000000000000"),
	(b"10000000001100100010011011101011", b"10000000000001100100101111101100"), -- 4.02749e-39 + -4.60574e-39 = -5.78249e-40
	(b"10000000000010000101110011000101", b"00000000000000000000000000000000"),
	(b"10000000010010101000001010110001", b"10000000010100101101111101110110"), -- -7.67963e-40 + -6.84271e-39 = -7.61067e-39
	(b"00000000011010010001110011110011", b"00000000000000000000000000000000"),
	(b"00000000000111011101100101010010", b"00000000100001101111011001000101"), -- 9.65311e-39 + 2.74119e-39 = 1.23943e-38
	(b"10000000000110111000000101011100", b"00000000000000000000000000000000"),
	(b"10000000001000001101000101101110", b"10000000001111000101001011001010"), -- -2.52596e-39 + -3.01387e-39 = -5.53983e-39
	(b"10000000001101001100110001011001", b"00000000000000000000000000000000"),
	(b"10000000011010100100100100010000", b"10000000100111110001010101101001"), -- -4.84875e-39 + -9.76077e-39 = -1.46095e-38
	(b"00000000010111011011110001001001", b"00000000000000000000000000000000"),
	(b"10000000010000100101111000111011", b"00000000000110110101111000001110"), -- 8.60825e-39 + -6.09495e-39 = 2.5133e-39
	(b"00000000000010011100101100100011", b"00000000000000000000000000000000"),
	(b"00000000001101010011001001011011", b"00000000001111101111110101111110"), -- 8.99391e-40 + 4.88535e-39 = 5.78474e-39
	(b"10000000000011101001100111101011", b"00000000000000000000000000000000"),
	(b"10000000001100111001010110101000", b"10000000010000100010111110010011"), -- -1.34091e-39 + -4.7373e-39 = -6.07821e-39
	(b"00000000010010101110101100100011", b"00000000000000000000000000000000"),
	(b"10000000001010010001110100101010", b"00000000001000011100110111111001"), -- 6.88018e-39 + -3.77572e-39 = 3.10446e-39
	(b"10000000000011000101010001011011", b"00000000000000000000000000000000"),
	(b"10000000011110100010001110111001", b"10000000100001100111100000010100"), -- -1.13229e-39 + -1.12167e-38 = -1.2349e-38
	(b"10000000001110000001001100100110", b"00000000000000000000000000000000"),
	(b"00000000001110000010000010000010", b"00000000000000000000110101011100"), -- -5.14966e-39 + 5.15445e-39 = 4.79244e-42
	(b"00000000010001011000111110000010", b"00000000000000000000000000000000"),
	(b"00000000000100001001001010001111", b"00000000010101100010001000010001"), -- 6.38813e-39 + 1.52194e-39 = 7.91007e-39
	(b"10000000011011110101000100000100", b"00000000000000000000000000000000"),
	(b"10000000011100110100100011010101", b"10000000111000101001100111011001"), -- -1.02228e-38 + -1.05872e-38 = -2.081e-38
	(b"00000000010100010110011011001111", b"00000000000000000000000000000000"),
	(b"10000000001010011000110011011011", b"00000000001001111101100111110100"), -- 7.47556e-39 + -3.81578e-39 = 3.65977e-39
	(b"10000000011100000000100000100111", b"00000000000000000000000000000000"),
	(b"10000000001010000101101001001101", b"10000000100110000110001001110100"), -- -1.02885e-38 + -3.70581e-39 = -1.39943e-38
	(b"00000000011110000110100100011101", b"00000000000000000000000000000000"),
	(b"10000000010101111011110001111101", b"00000000001000001010110010100000"), -- 1.1058e-38 + -8.05731e-39 = 3.00066e-39
	(b"00000000000001000100011110100101", b"00000000000000000000000000000000"),
	(b"00000000010100011010001100101111", b"00000000010101011110101011010100"), -- 3.93043e-40 + 7.49721e-39 = 7.89026e-39
	(b"10000000001011011000001101110011", b"00000000000000000000000000000000"),
	(b"00000000010100000110011111001111", b"00000000001000101110010001011100"), -- -4.17975e-39 + 7.38408e-39 = 3.20433e-39
	(b"00000000011001100000001110100011", b"00000000000000000000000000000000"),
	(b"10000000000011011111110011000011", b"00000000010110000000011011100000"), -- 9.36853e-39 + -1.28454e-39 = 8.08399e-39
	(b"10000000011101100011111100100011", b"00000000000000000000000000000000"),
	(b"10000000000111011100101111010101", b"10000000100101000000101011111000"), -- -1.08592e-38 + -2.73635e-39 = -1.35956e-38
	(b"00000000010110101011010111111110", b"00000000000000000000000000000000"),
	(b"00000000001000000111001111010011", b"00000000011110110010100111010001"), -- 8.33048e-39 + 2.98029e-39 = 1.13108e-38
	(b"00000000010011000101000011001100", b"00000000000000000000000000000000"),
	(b"00000000000101000010110000100011", b"00000000011000000111110011101111"), -- 7.00848e-39 + 1.85254e-39 = 8.86103e-39
	(b"10000000001011000111111111000100", b"00000000000000000000000000000000"),
	(b"10000000011010111010101111111000", b"10000000100110000010101110111100"), -- -4.0866e-39 + -9.88809e-39 = -1.39747e-38
	(b"00000000010111010011100110101100", b"00000000000000000000000000000000"),
	(b"10000000011011111011010101001000", b"10000000000100100111101110011100"), -- 8.56139e-39 + -1.02588e-38 = -1.69738e-39
	(b"00000000011111101001010001110110", b"00000000000000000000000000000000"),
	(b"10000000001001100110111011010101", b"00000000010110000010010110100001"), -- 1.16245e-38 + -3.52951e-39 = 8.09502e-39
	(b"00000000000111011111001110100100", b"00000000000000000000000000000000"),
	(b"10000000000000011101100110100011", b"00000000000111000001101000000001"), -- 2.75063e-39 + -1.69909e-40 = 2.58072e-39
	(b"10000000011001001001010001011011", b"00000000000000000000000000000000"),
	(b"10000000001001000000100000110101", b"10000000100010001001110010010000"), -- -9.23677e-39 + -3.30902e-39 = -1.25458e-38
	(b"00000000011111101001011000100000", b"00000000000000000000000000000000"),
	(b"00000000010110010000101011010100", b"00000000110101111010000011110100"), -- 1.16251e-38 + 8.17724e-39 = 1.98024e-38
	(b"10000000000010010000000110110100", b"00000000000000000000000000000000"),
	(b"00000000000011110110011010111110", b"00000000000001100110010100001010"), -- -8.2713e-40 + 1.41439e-39 = 5.87259e-40
	(b"00000000011111110101110100011101", b"00000000000000000000000000000000"),
	(b"10000000000000110010100111100110", b"00000000011111000011001100110111"), -- 1.16965e-38 + -2.90537e-40 = 1.1406e-38
	(b"10000000011000100111111101111100", b"00000000000000000000000000000000"),
	(b"00000000010001000010111010111000", b"10000000000111100101000011000100"), -- -9.04561e-39 + 6.26157e-39 = -2.78404e-39
	(b"10000000001110010011011110011011", b"00000000000000000000000000000000"),
	(b"10000000000011100000000000000111", b"10000000010001110011011110100010"), -- -5.25457e-39 + -1.28571e-39 = -6.54028e-39
	(b"00000000000111110011110111000101", b"00000000000000000000000000000000"),
	(b"10000000001010001010001011111100", b"10000000000010010110010100110111"), -- 2.86906e-39 + -3.73189e-39 = -8.62829e-40
	(b"00000000000001000010010001110000", b"00000000000000000000000000000000"),
	(b"10000000011001110010010111110001", b"10000000011000110000000110000001"), -- 3.80413e-40 + -9.47267e-39 = -9.09225e-39
	(b"00000000010001010101110010000101", b"00000000000000000000000000000000"),
	(b"10000000011000000001100010010101", b"10000000000110101011110000010000"), -- 6.36984e-39 + -8.82503e-39 = -2.45519e-39
	(b"10000000000101101000011011111010", b"00000000000000000000000000000000"),
	(b"10000000000101000011100000011100", b"10000000001010101011111100010110"), -- -2.0688e-39 + -1.85684e-39 = -3.92564e-39
	(b"10000000011110111011111000101110", b"00000000000000000000000000000000"),
	(b"10000000010001000000100101110011", b"10000000101111111100011110100001"), -- -1.1364e-38 + -6.2482e-39 = -1.76122e-38
	(b"10000000000101010001000001111011", b"00000000000000000000000000000000"),
	(b"00000000001011101010110101001111", b"00000000000110011001110011010100"), -- -1.93446e-39 + 4.2866e-39 = 2.35215e-39
	(b"00000000001110100100100010100010", b"00000000000000000000000000000000"),
	(b"00000000001111110010111010100011", b"00000000011110010111011101000101"), -- 5.35251e-39 + 5.80237e-39 = 1.11549e-38
	(b"00000000001111001101011100101010", b"00000000000000000000000000000000"),
	(b"00000000010110011001101111111011", b"00000000100101100111001100100101"), -- 5.58732e-39 + 8.22931e-39 = 1.38166e-38
	(b"00000000011010100010110010101101", b"00000000000000000000000000000000"),
	(b"00000000000010001000111110110011", b"00000000011100101011110001100000"), -- 9.75059e-39 + 7.86234e-40 = 1.05368e-38
	(b"00000000001111000010101101101100", b"00000000000000000000000000000000"),
	(b"10000000001010010110100010010011", b"00000000000100101100001011011001"), -- 5.52571e-39 + -3.80277e-39 = 1.72294e-39
	(b"10000000011000001101010010100110", b"00000000000000000000000000000000"),
	(b"10000000000011101110101110101010", b"10000000011011111100000001010000"), -- -8.89249e-39 + -1.37024e-39 = -1.02627e-38
	(b"00000000010010011100111111101000", b"00000000000000000000000000000000"),
	(b"00000000010000001100011000100100", b"00000000100010101001011000001100"), -- 6.77857e-39 + 5.94855e-39 = 1.27271e-38
	(b"00000000001110001000100001110101", b"00000000000000000000000000000000"),
	(b"00000000011101101010101100111111", b"00000000101011110011001110110100"), -- 5.19174e-39 + 1.0898e-38 = 1.60898e-38
	(b"10000000000010110000100001101101", b"00000000000000000000000000000000"),
	(b"00000000011010111101000000010001", b"00000000011000001100011110100100"), -- -1.01321e-39 + 9.90104e-39 = 8.88783e-39
	(b"10000000011110111110000000010001", b"00000000000000000000000000000000"),
	(b"00000000011001011001111001000000", b"10000000000101100100000111010001"), -- -1.13761e-38 + 9.33215e-39 = -2.04399e-39
	(b"10000000000101001100001101101101", b"00000000000000000000000000000000"),
	(b"00000000001100100110010110010111", b"00000000000111011010001000101010"), -- -1.90682e-39 + 4.62822e-39 = 2.7214e-39
	(b"00000000011101111111111100011010", b"00000000000000000000000000000000"),
	(b"00000000001111010001100111010000", b"00000000101101010001100011101010"), -- 1.10199e-38 + 5.61123e-39 = 1.66312e-38
	(b"00000000001000100001010100011010", b"00000000000000000000000000000000"),
	(b"00000000001111011111000100100011", b"00000000011000000000011000111101"), -- 3.12998e-39 + 5.68847e-39 = 8.81845e-39
	(b"10000000001110101101100100010100", b"00000000000000000000000000000000"),
	(b"10000000010011100101111010101111", b"10000000100010010011011111000011"), -- -5.40433e-39 + -7.19713e-39 = -1.26015e-38
	(b"10000000001101110001010100110100", b"00000000000000000000000000000000"),
	(b"10000000001101101001110100110111", b"10000000011011011011001001101011"), -- -5.05856e-39 + -5.01551e-39 = -1.00741e-38
	(b"10000000000011111110111001010101", b"00000000000000000000000000000000"),
	(b"00000000000101001111110111100001", b"00000000000001010000111110001100"), -- -1.46303e-39 + 1.92778e-39 = 4.64755e-40
	(b"10000000010010110000000011000000", b"00000000000000000000000000000000"),
	(b"10000000010100101101100100100011", b"10000000100111011101100111100011"), -- -6.88793e-39 + -7.6084e-39 = -1.44963e-38
	(b"00000000000011010001010111010110", b"00000000000000000000000000000000"),
	(b"10000000000011100101111011110110", b"10000000000000010100100100100000"), -- 1.20169e-39 + -1.31976e-39 = -1.18068e-40
	(b"00000000011001011100001011110001", b"00000000000000000000000000000000"),
	(b"10000000011010010110100010111100", b"10000000000000111010010111001011"), -- 9.34532e-39 + -9.6803e-39 = -3.34982e-40
	(b"10000000010111110011001010010001", b"00000000000000000000000000000000"),
	(b"00000000010110100100101001111000", b"10000000000001001110100000011001"), -- -8.74251e-39 + 8.29191e-39 = -4.50603e-40
	(b"10000000001011010110010111010111", b"00000000000000000000000000000000"),
	(b"00000000000001110101001010011010", b"10000000001001100001001100111101"), -- -4.16913e-39 + 6.7248e-40 = -3.49665e-39
	(b"00000000001001000101110101011011", b"00000000000000000000000000000000"),
	(b"00000000000110101100010000000111", b"00000000001111110010000101100010"), -- 3.33957e-39 + 2.45804e-39 = 5.79761e-39
	(b"10000000011000000110001110011100", b"00000000000000000000000000000000"),
	(b"00000000000000111011010110110001", b"10000000010111001010110111101011"), -- -8.85194e-39 + 3.40685e-40 = -8.51126e-39
	(b"00000000001111011110010000001011", b"00000000000000000000000000000000"),
	(b"00000000001001011001110000001110", b"00000000011000111000000000011001"), -- 5.68377e-39 + 3.4539e-39 = 9.13767e-39
	(b"10000000001100000011011001011010", b"00000000000000000000000000000000"),
	(b"10000000001110001100110001001100", b"10000000011010010000001010100110"), -- -4.4276e-39 + -5.21608e-39 = -9.64368e-39
	(b"00000000001110000101001100111111", b"00000000000000000000000000000000"),
	(b"00000000011101100100001100001101", b"00000000101011101001011001001100"), -- 5.17265e-39 + 1.08606e-38 = 1.60333e-38
	(b"10000000011101011011100101110111", b"00000000000000000000000000000000"),
	(b"10000000011000000001001011100001", b"10000000110101011100110001011000"), -- -1.08113e-38 + -8.82298e-39 = -1.96343e-38
	(b"00000000001101011110110110000101", b"00000000000000000000000000000000"),
	(b"10000000011011011111111101101000", b"10000000001110000001000111100011"), -- 4.95249e-39 + -1.01017e-38 = -5.1492e-39
	(b"10000000000110111110001100000110", b"00000000000000000000000000000000"),
	(b"00000000001101111110000101111110", b"00000000000110111111111001111000"), -- -2.561e-39 + 5.13184e-39 = 2.57084e-39
	(b"00000000010111100011011000011111", b"00000000000000000000000000000000"),
	(b"00000000011111011110100000010000", b"00000000110111000001111000101111"), -- 8.65195e-39 + 1.15627e-38 = 2.02146e-38
	(b"10000000011011110110000000011011", b"00000000000000000000000000000000"),
	(b"10000000011101100100011101110000", b"10000000111001011010011110001011"), -- -1.02282e-38 + -1.08622e-38 = -2.10904e-38
	(b"10000000001110101100111101110001", b"00000000000000000000000000000000"),
	(b"10000000010011100100101000100101", b"10000000100010010001100110010110"), -- -5.40087e-39 + -7.18977e-39 = -1.25906e-38
	(b"10000000001011011100010000110100", b"00000000000000000000000000000000"),
	(b"00000000000011000011000111011111", b"10000000001000011001001001010101"), -- -4.20298e-39 + 1.11992e-39 = -3.08307e-39
	(b"00000000000101000011011011000100", b"00000000000000000000000000000000"),
	(b"10000000011011110100111110001110", b"10000000010110110001100011001010"), -- 1.85636e-39 + -1.02223e-38 = -8.36592e-39
	(b"10000000011110100000110001110101", b"00000000000000000000000000000000"),
	(b"00000000011100001110000001001001", b"10000000000010010010110000101100"), -- -1.12084e-38 + 1.0366e-38 = -8.42365e-40
	(b"00000000010001100110101000101111", b"00000000000000000000000000000000"),
	(b"00000000001110010010000110011110", b"00000000011111111000101111001101"), -- 6.46658e-39 + 5.24668e-39 = 1.17133e-38
	(b"10000000010110010111110000001000", b"00000000000000000000000000000000"),
	(b"00000000000010101111011011000110", b"10000000010011101000010101000010"), -- -8.21785e-39 + 1.00688e-39 = -7.21097e-39
	(b"00000000010000101101110101100010", b"00000000000000000000000000000000"),
	(b"00000000000011000110101010001111", b"00000000010011110100011111110001"), -- 6.14056e-39 + 1.14025e-39 = 7.28081e-39
	(b"10000000000101000000101110111000", b"00000000000000000000000000000000"),
	(b"10000000010111010101011111000010", b"10000000011100010110001101111010"), -- -1.84091e-39 + -8.57218e-39 = -1.04131e-38
	(b"00000000000111100010010111001001", b"00000000000000000000000000000000"),
	(b"00000000001111101111101110100101", b"00000000010111010010000101101110"), -- 2.76862e-39 + 5.78407e-39 = 8.55269e-39
	(b"10000000010100101011000000010100", b"00000000000000000000000000000000"),
	(b"00000000000000101001011011110100", b"10000000010100000001100100100000"), -- -7.59368e-39 + 2.37823e-40 = -7.35585e-39
	(b"00000000000110111010011101101000", b"00000000000000000000000000000000"),
	(b"00000000001100100101111001001001", b"00000000010011100000010110110001"), -- 2.53961e-39 + 4.6256e-39 = 7.16521e-39
	(b"10000000000101111111011001011010", b"00000000000000000000000000000000"),
	(b"10000000001000010011001101001101", b"10000000001110010010100110100111"), -- -2.20059e-39 + -3.04897e-39 = -5.24957e-39
	(b"00000000010011110110101011101110", b"00000000000000000000000000000000"),
	(b"00000000001011001101111101101101", b"00000000011111000100101001011011"), -- 7.29336e-39 + 4.12091e-39 = 1.14143e-38
	(b"00000000011010110001110110011001", b"00000000000000000000000000000000"),
	(b"10000000011111010011011101001100", b"10000000000100100001100110110011"), -- 9.83702e-39 + -1.14993e-38 = -1.66226e-39
	(b"10000000000110100110001111000010", b"00000000000000000000000000000000"),
	(b"00000000011001111101001101000101", b"00000000010011010110111110000011"), -- -2.42351e-39 + 9.53485e-39 = 7.11134e-39
	(b"10000000000100010011100111000000", b"00000000000000000000000000000000"),
	(b"00000000001001101101010111101001", b"00000000000101011001110000101001"), -- -1.58192e-39 + 3.56649e-39 = 1.98457e-39
	(b"10000000010100000101001010101110", b"00000000000000000000000000000000"),
	(b"10000000001010111100100110111001", b"10000000011111000001110001100111"), -- -7.3765e-39 + -4.02129e-39 = -1.13978e-38
	(b"10000000010000010011010110001100", b"00000000000000000000000000000000"),
	(b"00000000011111001011001011011010", b"00000000001110110111110101001110"), -- -5.98852e-39 + 1.14518e-38 = 5.46325e-39
	(b"00000000001001001011100000100010", b"00000000000000000000000000000000"),
	(b"00000000010111110101011101011110", b"00000000100001000000111110000000"), -- 3.37213e-39 + 8.75571e-39 = 1.21278e-38
	(b"00000000000000101101100011111110", b"00000000000000000000000000000000"),
	(b"10000000001110111101000101101001", b"10000000001110001111100001101011"), -- 2.61513e-40 + -5.49342e-39 = -5.2319e-39
	(b"10000000011110000110101101010100", b"00000000000000000000000000000000"),
	(b"10000000000100101101011110000001", b"10000000100010110100001011010101"), -- -1.10588e-38 + -1.73035e-39 = -1.27891e-38
	(b"00000000010001011100100111111101", b"00000000000000000000000000000000"),
	(b"00000000000010010100001000110100", b"00000000010011110000110000110001"), -- 6.40911e-39 + 8.50269e-40 = 7.25938e-39
	(b"00000000001000001011111010100010", b"00000000000000000000000000000000"),
	(b"10000000000000000110100001010001", b"00000000001000000101011001010001"), -- 3.00712e-39 + -3.74217e-41 = 2.9697e-39
	(b"10000000011011000101110110110100", b"00000000000000000000000000000000"),
	(b"00000000001011000000101001101000", b"10000000010000000101001101001100"), -- -9.95185e-39 + 4.04449e-39 = -5.90735e-39
	(b"00000000011110000001111101111010", b"00000000000000000000000000000000"),
	(b"10000000001000111111010111010000", b"00000000010101000010100110101010"), -- 1.10316e-38 + -3.30242e-39 = 7.72913e-39
	(b"00000000010010100110111010101011", b"00000000000000000000000000000000"),
	(b"10000000011011010010100101101001", b"10000000001000101011101010111110"), -- 6.83553e-39 + -1.00249e-38 = -3.1894e-39
	(b"00000000001111010100111101110110", b"00000000000000000000000000000000"),
	(b"00000000010111101011111111110110", b"00000000100111000000111101101100"), -- 5.63047e-39 + 8.7014e-39 = 1.43319e-38
	(b"01110000001101000011111011110001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.23134e+29 + inf = inf
	(b"10100001101000110000000000101010", b"00000000000000000000000000000000"),
	(b"10010000100101010011010101111100", b"10100001101000110000000000101010"), -- -1.10454e-18 + -5.88525e-29 = -1.10454e-18
	(b"10100101111010110110111100010000", b"00000000000000000000000000000000"),
	(b"10100110111010100111100100101000", b"10100111000100101010101001110110"), -- -4.08413e-16 + -1.62699e-15 = -2.0354e-15
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100110000101001010001011100010", b"11100110000101001010001011100010"), -- -0 + -1.75479e+23 = -1.75479e+23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110010110100010011110000001010", b"00110010110100010011110000001010"), -- 0 + 2.43581e-08 = 2.43581e-08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010100110110000110111001101001", b"01111111100000000000000000000000"), -- inf + 7.43652e+12 = inf
	(b"11011100110000011010101110101011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000011", b"11011100110000011010101110101011"), -- -4.36107e+17 + -4.2039e-45 = -4.36107e+17
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11110100011111010111111010111100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110100011111010111111010111100"), -- -8.03358e+31 + -0 = -8.03358e+31
	(b"11001000010000010100101010000110", b"00000000000000000000000000000000"),
	(b"11011101111011100101111000000110", b"11011101111011100101111000000110"), -- -197930 + -2.14702e+18 = -2.14702e+18
	(b"00010000000001000010100101100111", b"00000000000000000000000000000000"),
	(b"00000111010110100010011010111011", b"00010000000001000010100110011110"), -- 2.60643e-29 + 1.64119e-34 = 2.60645e-29
	(b"00100100111011010011010001000010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.02871e-16 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100000000001111000110101010110", b"10100000000001111000110101010110"), -- -0 + -1.14817e-19 = -1.14817e-19
	(b"10001110111101110100011100000011", b"00000000000000000000000000000000"),
	(b"11010111111110100111100100101000", b"11010111111110100111100100101000"), -- -6.09586e-30 + -5.50797e+14 = -5.50797e+14
	(b"01000111010110001110010011010001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 55524.8 + inf = inf
	(b"01010011101010011100100101111011", b"00000000000000000000000000000000"),
	(b"01100000100000100000000000111111", b"01100000100000100000000000111111"), -- 1.45846e+12 + 7.49405e+19 = 7.49405e+19
	(b"11100011011011101110101000001111", b"00000000000000000000000000000000"),
	(b"11110100100110001001011111010010", b"11110100100110001001011111010010"), -- -4.40719e+21 + -9.67173e+31 = -9.67173e+31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111101100111111001101000111001", b"11111111100000000000000000000000"), -- -inf + -2.65185e+37 = -inf
	(b"01101010000100101011000000111110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.43339e+25 + inf = inf
	(b"01100001010100001011001010100010", b"00000000000000000000000000000000"),
	(b"01110110011001001101111010000001", b"01110110011001001101111010000001"), -- 2.40612e+20 + 1.1605e+33 = 1.1605e+33
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00110010011111111101010110110011", b"00000000000000000000000000000000"),
	(b"00100001000111101111011010100001", b"00110010011111111101010110110011"), -- 1.48915e-08 + 5.38589e-19 = 1.48915e-08
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001000100100110000100101101110", b"01001000100100110000100101101110"), -- 0 + 301131 = 301131
	(b"11001011111010111101100101000110", b"00000000000000000000000000000000"),
	(b"10111001010001011110011100000101", b"11001011111010111101100101000110"), -- -3.09132e+07 + -0.000188734 = -3.09132e+07
	(b"11101111100110100010010111100010", b"00000000000000000000000000000000"),
	(b"10110001101010101010101110111010", b"11101111100110100010010111100010"), -- -9.5413e+28 + -4.96717e-09 = -9.5413e+28
	(b"01110111101001000101101111101011", b"00000000000000000000000000000000"),
	(b"01101000000110101010001011110111", b"01110111101001000101101111101011"), -- 6.6672e+33 + 2.921e+24 = 6.6672e+33
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001000101011010100110111000101", b"01111111100000000000000000000000"), -- inf + 354926 = inf
	(b"11101011101010100001001101101010", b"00000000000000000000000000000000"),
	(b"11001110100110000000001100101000", b"11101011101010100001001101101010"), -- -4.11218e+26 + -1.27517e+09 = -4.11218e+26
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010000111011000000000010111011", b"11111111100000000000000000000000"), -- -inf + -3.16758e+10 = -inf
	(b"10000000000000000000000101111011", b"00000000000000000000000000000000"),
	(b"11010000100101001100100010010110", b"11010000100101001100100010010110"), -- -5.31092e-43 + -1.99694e+10 = -1.99694e+10
	(b"01010010100111111111011111001101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.43529e+11 + inf = inf
	(b"00011011001000111000110001110101", b"00000000000000000000000000000000"),
	(b"00100110000000010000101000110111", b"00100110000000010000101000111010"), -- 1.35284e-22 + 4.47697e-16 = 4.47697e-16
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111001111111010101011111111101", b"10111001111111010101011111111101"), -- -0 + -0.000483215 = -0.000483215
	(b"10000000000001101010010101110011", b"00000000000000000000000000000000"),
	(b"11011101001011110100110110100010", b"11011101001011110100110110100010"), -- -6.10365e-40 + -7.89496e+17 = -7.89496e+17
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001100111101101110110110011011", b"11111111100000000000000000000000"), -- -inf + -3.80453e-31 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010001000000111101111010001000", b"11111111100000000000000000000000"), -- -inf + -1.04027e-28 = -inf
	(b"01010011011111001001011010100000", b"00000000000000000000000000000000"),
	(b"01010011110101110111110000001010", b"01010100001010101110001110101101"), -- 1.08486e+12 + 1.851e+12 = 2.93586e+12
	(b"11001101101110010101011110001110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.8869e+08 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000111100110011000000110100101", b"11111111100000000000000000000000"), -- -inf + -78595.3 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100010011110001101000111110011", b"11111111100000000000000000000000"), -- -inf + -3.37214e-18 = -inf
	(b"11001110100110100011001111000100", b"00000000000000000000000000000000"),
	(b"11001001101110001100101001111111", b"11001110100110100110000111110111"), -- -1.29354e+09 + -1.51381e+06 = -1.29506e+09
	(b"00111100100010001001011111111100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000001101011", b"00111100100010001001011111111100"), -- 0.016674 + 1.49939e-43 = 0.016674
	(b"10010000101011001111101110000000", b"00000000000000000000000000000000"),
	(b"11010000000000011101101001011011", b"11010000000000011101101001011011"), -- -6.82295e-29 + -8.71428e+09 = -8.71428e+09
	(b"00000000000001011100100110010011", b"00000000000000000000000000000000"),
	(b"00100110000111011000000111001100", b"00100110000111011000000111001100"), -- 5.31489e-40 + 5.46462e-16 = 5.46462e-16
	(b"10100100100011001101000001101000", b"00000000000000000000000000000000"),
	(b"10101010100111001111011110011111", b"10101010100111010000000001101100"), -- -6.10684e-17 + -2.7883e-13 = -2.78891e-13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001101011110100000010011001101", b"01111111100000000000000000000000"), -- inf + 2.62164e+08 = inf
	(b"01011000101010110010000001011001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.50524e+15 + inf = inf
	(b"01111001100000111111100011000111", b"00000000000000000000000000000000"),
	(b"01001100111110011010001000110100", b"01111001100000111111100011000111"), -- 8.56546e+34 + 1.3088e+08 = 8.56546e+34
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110010111110001000110011000101", b"00110010111110001000110011000101"), -- 0 + 2.8935e-08 = 2.8935e-08
	(b"11111101011000111011011111110010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.89181e+37 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00111101001010010001000100111011", b"00000000000000000000000000000000"),
	(b"01111110100101101100100000111111", b"01111110100101101100100000111111"), -- 0.0412762 + 1.00212e+38 = 1.00212e+38
	(b"01111110011111011011010001011011", b"00000000000000000000000000000000"),
	(b"00010111001010000101011000100101", b"01111110011111011011010001011011"), -- 8.43078e+37 + 5.43925e-25 = 8.43078e+37
	(b"00101101001001001001000000101010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.35433e-12 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001100001101110110001010110100", b"01001100001101110110001010110100"), -- 0 + 4.80734e+07 = 4.80734e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010011000001110011100011100100", b"11010011000001110011100011100100"), -- -0 + -5.80775e+11 = -5.80775e+11
	(b"11110001110001100000010010010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.96107e+30 + -inf = -inf
	(b"01010110100010111011000010111000", b"00000000000000000000000000000000"),
	(b"01111111001111100010011000010110", b"01111111001111100010011000010110"), -- 7.67956e+13 + 2.52751e+38 = 2.52751e+38
	(b"11001110000011000011001001000010", b"00000000000000000000000000000000"),
	(b"11011010101100001011001100011101", b"11011010101100001011001100011101"), -- -5.88026e+08 + -2.48683e+16 = -2.48683e+16
	(b"10000000001100110011101110010001", b"00000000000000000000000000000000"),
	(b"11001101010001001100101000001001", b"11001101010001001100101000001001"), -- -4.70498e-39 + -2.06348e+08 = -2.06348e+08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100010011000011010000001001110", b"01111111100000000000000000000000"), -- inf + 1.04052e+21 = inf
	(b"00111101101010101110101010011100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111101101010101110101010011100"), -- 0.0834553 + 0 = 0.0834553
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001001010000001111010011010111", b"10001001010000001111010011010111"), -- -0 + -2.32263e-33 = -2.32263e-33
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000001001110001010001", b"00000000000000000000000000000000"),
	(b"10011101000100111110111001101000", b"10011101000100111110111001101000"), -- -5.60758e-41 + -1.95785e-21 = -1.95785e-21
	(b"01000100111111111010101100011110", b"00000000000000000000000000000000"),
	(b"00000001101010100111110110111110", b"01000100111111111010101100011110"), -- 2045.35 + 6.26286e-38 = 2045.35
	(b"00011100000010101010101101010100", b"00000000000000000000000000000000"),
	(b"01101101000111011100111011101000", b"01101101000111011100111011101000"), -- 4.58818e-22 + 3.05246e+27 = 3.05246e+27
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110110010100010100110010000100", b"11111111100000000000000000000000"), -- -inf + -3.1188e-06 = -inf
	(b"11100111101100101100001111010110", b"00000000000000000000000000000000"),
	(b"10010011100001000101111000000101", b"11100111101100101100001111010110"), -- -1.68839e+24 + -3.34142e-27 = -1.68839e+24
	(b"00000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000001"), -- 1.4013e-45 + 0 = 1.4013e-45
	(b"11000011000110101111100011100011", b"00000000000000000000000000000000"),
	(b"10111110101001100110001010011001", b"11000011000110110100110000010100"), -- -154.972 + -0.324971 = -155.297
	(b"00100000110100010011001000111010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.54392e-19 + inf = inf
	(b"00110110010110001011000111100101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00110110010110001011000111100101"), -- 3.22901e-06 + 0 = 3.22901e-06
	(b"01010101101001011000100010010001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.27507e+13 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000010011101000111101011010111", b"01111111100000000000000000000000"), -- inf + 1.79615e-37 = inf
	(b"00101011100111111110000001101001", b"00000000000000000000000000000000"),
	(b"01011011110110100000001110000111", b"01011011110110100000001110000111"), -- 1.13599e-12 + 1.22731e+17 = 1.22731e+17
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001011011101101000100110111", b"11111111100000000000000000000000"), -- -inf + -1.80445e+25 = -inf
	(b"00111111100110110101001011011000", b"00000000000000000000000000000000"),
	(b"01000111000100100000000110101010", b"01000111000100100000001011100001"), -- 1.21347 + 37377.7 = 37378.9
	(b"10010011110011100000000101011111", b"00000000000000000000000000000000"),
	(b"11000101010010011110001001010001", b"11000101010010011110001001010001"), -- -5.20031e-27 + -3230.14 = -3230.14
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001010110110101100001100110000", b"00001010110110101100001100110000"), -- 0 + 2.10661e-32 = 2.10661e-32
	(b"11101110001001101100110110001011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.29057e+28 + -inf = -inf
	(b"11101111001000010001011011011101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11101111001000010001011011011101"), -- -4.98547e+28 + -0 = -4.98547e+28
	(b"00110011111100101111110000100101", b"00000000000000000000000000000000"),
	(b"01100111010001001000000101011011", b"01100111010001001000000101011011"), -- 1.13149e-07 + 9.2797e+23 = 9.2797e+23
	(b"01001001010010100111111110101111", b"00000000000000000000000000000000"),
	(b"00101111100110110111011000000011", b"01001001010010100111111110101111"), -- 829435 + 2.82782e-10 = 829435
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00001011100111110101011010001010", b"00000000000000000000000000000000"),
	(b"01110111001011001101111101010110", b"01110111001011001101111101010110"), -- 6.13748e-32 + 3.50627e+33 = 3.50627e+33
	(b"10101101010000001001001111111110", b"00000000000000000000000000000000"),
	(b"11100111010111110001001000101010", b"11100111010111110001001000101010"), -- -1.09468e-11 + -1.05342e+24 = -1.05342e+24
	(b"00101110001100011010100111101001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00101110001100011010100111101001"), -- 4.03961e-11 + 0 = 4.03961e-11
	(b"10111011000101010011000101111100", b"00000000000000000000000000000000"),
	(b"10101100100110111011000111111100", b"10111011000101010011000101111100"), -- -0.00227651 + -4.42513e-12 = -0.00227651
	(b"11100110100100001000011001111111", b"00000000000000000000000000000000"),
	(b"11001100010011100010011101010111", b"11100110100100001000011001111111"), -- -3.41251e+23 + -5.40419e+07 = -3.41251e+23
	(b"11001000001001001110011000001000", b"00000000000000000000000000000000"),
	(b"11010011011010001011101011000001", b"11010011011010001011101011000100"), -- -168856 + -9.99566e+11 = -9.99566e+11
	(b"00101110010111000111010100111101", b"00000000000000000000000000000000"),
	(b"00010110110001100100101000010101", b"00101110010111000111010100111101"), -- 5.01263e-11 + 3.20354e-25 = 5.01263e-11
	(b"01110100101101000000011000001110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01110100101101000000011000001110"), -- 1.14104e+32 + 0 = 1.14104e+32
	(b"10111011100101011110101110111101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0.00457522 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100010010011001111110111101010", b"00100010010011001111110111101010"), -- 0 + 2.77816e-18 = 2.77816e-18
	(b"00101101000110011100111001111101", b"00000000000000000000000000000000"),
	(b"01111011011000001000000110001010", b"01111011011000001000000110001010"), -- 8.74289e-12 + 1.1657e+36 = 1.1657e+36
	(b"10100001010111000001000000110010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.45603e-19 + -inf = -inf
	(b"10000000000000001101111101101011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.01473e-41 + -inf = -inf
	(b"10010010000000100100011001100000", b"00000000000000000000000000000000"),
	(b"10110000100001101110010001110101", b"10110000100001101110010001110101"), -- -4.11075e-28 + -9.81471e-10 = -9.81471e-10
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000001001111111", b"10000000000000000000001001111111"), -- -0 + -8.9543e-43 = -8.9543e-43
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01000010011011101010101111011000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 59.6678 + inf = inf
	(b"11110111101001110011001111001000", b"00000000000000000000000000000000"),
	(b"10000100111110000100100011010101", b"11110111101001110011001111001000"), -- -6.78253e+33 + -5.83714e-36 = -6.78253e+33
	(b"00110011111110101011111101010100", b"00000000000000000000000000000000"),
	(b"01101100100101001001100101010011", b"01101100100101001001100101010011"), -- 1.16763e-07 + 1.43716e+27 = 1.43716e+27
	(b"11011010101111101110110000100000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.68699e+16 + -inf = -inf
	(b"10000000000000000000000000011010", b"00000000000000000000000000000000"),
	(b"10000110100001111011110110110011", b"10000110100001111011110110110011"), -- -3.64338e-44 + -5.10601e-35 = -5.10601e-35
	(b"01110101000111110000010111011100", b"00000000000000000000000000000000"),
	(b"00100000000000100101011100011100", b"01110101000111110000010111011100"), -- 2.01585e+32 + 1.10403e-19 = 2.01585e+32
	(b"01111101011101010001010001000110", b"00000000000000000000000000000000"),
	(b"01010111100011100101110100110110", b"01111101011101010001010001000110"), -- 2.03604e+37 + 3.13062e+14 = 2.03604e+37
	(b"10001101010111011010110010010111", b"00000000000000000000000000000000"),
	(b"10011111000111100111000001010110", b"10011111000111100111000001010110"), -- -6.83086e-31 + -3.35507e-20 = -3.35507e-20
	(b"10000110110100111100101111101110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.9669e-35 + -inf = -inf
	(b"10001000101101110100000110000001", b"00000000000000000000000000000000"),
	(b"11000011100100100100011101100110", b"11000011100100100100011101100110"), -- -1.10293e-33 + -292.558 = -292.558
	(b"00110011101110111010110101010010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 8.73939e-08 + inf = inf
	(b"00110011011100111100001100111001", b"00000000000000000000000000000000"),
	(b"01001001100010101110100110000111", b"01001001100010101110100110000111"), -- 5.67554e-08 + 1.13797e+06 = 1.13797e+06
	(b"10011111000000001110110001000100", b"00000000000000000000000000000000"),
	(b"11010010101011000110100011110100", b"11010010101011000110100011110100"), -- -2.73005e-20 + -3.70248e+11 = -3.70248e+11
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010111001000010011100000010001", b"11111111100000000000000000000000"), -- -inf + -1.77262e+14 = -inf
	(b"11000110100101101101000011101101", b"00000000000000000000000000000000"),
	(b"11011101010011001100010101000001", b"11011101010011001100010101000001"), -- -19304.5 + -9.22204e+17 = -9.22204e+17
	(b"10100101101010110011010000011011", b"00000000000000000000000000000000"),
	(b"10011110111101010110100100111110", b"10100101101010110011011111110001"), -- -2.96991e-16 + -2.59839e-20 = -2.97017e-16
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000010110", b"10000000000000000000000000010110"), -- -0 + -3.08286e-44 = -3.08286e-44
	(b"00101011001000001001101110110100", b"00000000000000000000000000000000"),
	(b"00101110101101110010111001011110", b"00101110101110000110111110010101"), -- 5.70595e-13 + 8.33011e-11 = 8.38717e-11
	(b"11100011000011100000001011011111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.61964e+21 + -inf = -inf
	(b"01010111100000000000001000100001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.81493e+14 + inf = inf
	(b"11000000001010000010010000100101", b"00000000000000000000000000000000"),
	(b"11101000101010011000111111110010", b"11101000101010011000111111110010"), -- -2.62721 + -6.40588e+24 = -6.40588e+24
	(b"11010101100000001110101000000110", b"00000000000000000000000000000000"),
	(b"11101101111001010110110101011011", b"11101101111001010110110101011011"), -- -1.77178e+13 + -8.87553e+27 = -8.87553e+27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010101100000101010111011011", b"11011010101100000101010111011011"), -- -0 + -2.4817e+16 = -2.4817e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001101000010111110100", b"11111111100000000000000000000000"), -- -inf + -2.60193 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000110111100011101011001011111", b"01111111100000000000000000000000"), -- inf + 30955.2 = inf
	(b"11000110110010011101110101010000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000110110010011101110101010000"), -- -25838.7 + -0 = -25838.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11010000101001100001010001101101", b"00000000000000000000000000000000"),
	(b"11000001010001100101111001001111", b"11010000101001100001010001101101"), -- -2.22909e+10 + -12.398 = -2.22909e+10
	(b"11101001001100111000000011101100", b"00000000000000000000000000000000"),
	(b"10001110010001011100101111011101", b"11101001001100111000000011101100"), -- -1.35629e+25 + -2.43803e-30 = -1.35629e+25
	(b"10001001011001011010111100011010", b"00000000000000000000000000000000"),
	(b"11000010100100100101010010111110", b"11000010100100100101010010111110"), -- -2.76472e-33 + -73.1655 = -73.1655
	(b"10101011110001111010100011110111", b"00000000000000000000000000000000"),
	(b"11000111110110001011111000100110", b"11000111110110001011111000100110"), -- -1.41867e-12 + -110972 = -110972
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110010011011011001101100101111", b"11111111100000000000000000000000"), -- -inf + -4.70628e+30 = -inf
	(b"01000111110001011011001001110101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000111110001011011001001110101"), -- 101221 + 0 = 101221
	(b"11010111000101100110100010111101", b"00000000000000000000000000000000"),
	(b"11100010100001100101110101001111", b"11100010100001100101110101010000"), -- -1.65377e+14 + -1.23929e+21 = -1.23929e+21
	(b"01111101010110101001010001000010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.81588e+37 + inf = inf
	(b"11101001010100101100110000011011", b"00000000000000000000000000000000"),
	(b"10001010100000010100010011010000", b"11101001010100101100110000011011"), -- -1.59274e+25 + -1.24481e-32 = -1.59274e+25
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100101100011111101011101001101", b"01111111100000000000000000000000"), -- inf + 8.49088e+22 = inf
	(b"11001000101010001010000100010100", b"00000000000000000000000000000000"),
	(b"11110001101101101000100111000111", b"11110001101101101000100111000111"), -- -345353 + -1.80777e+30 = -1.80777e+30
	(b"00000000000000000000100110101010", b"00000000000000000000000000000000"),
	(b"01001011010100010001010101011100", b"01001011010100010001010101011100"), -- 3.46681e-42 + 1.37025e+07 = 1.37025e+07
	(b"00100001110001010001111101011011", b"00000000000000000000000000000000"),
	(b"01110010000001100011110111000001", b"01110010000001100011110111000001"), -- 1.33575e-18 + 2.65892e+30 = 2.65892e+30
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001100100001010110111010101100", b"01111111100000000000000000000000"), -- inf + 6.9957e+07 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001001000001100000101010000111", b"11111111100000000000000000000000"), -- -inf + -549032 = -inf
	(b"00000000000000000001111101111100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.12945e-41 + inf = inf
	(b"01111001110010111101001011111011", b"00000000000000000000000000000000"),
	(b"01011110000100100101010110001000", b"01111001110010111101001011111011"), -- 1.32289e+35 + 2.63612e+18 = 1.32289e+35
	(b"00100110100010110010111010001010", b"00000000000000000000000000000000"),
	(b"00110111011010100001111110101011", b"00110111011010100001111110101011"), -- 9.65768e-16 + 1.39549e-05 = 1.39549e-05
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101000101100000101010101010100", b"11111111100000000000000000000000"), -- -inf + -1.95769e-14 = -inf
	(b"10011101000110111100010100111101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.0616e-21 + -inf = -inf
	(b"10100001110100010111111011110001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.4196e-18 + -inf = -inf
	(b"10010110011101100000110100111011", b"00000000000000000000000000000000"),
	(b"11001111101011100000111110000010", b"11001111101011100000111110000010"), -- -1.98759e-25 + -5.8405e+09 = -5.8405e+09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110110011000000000111100100111", b"01111111100000000000000000000000"), -- inf + 1.13612e+33 = inf
	(b"00111010001001111001110101010111", b"00000000000000000000000000000000"),
	(b"00011010111100000011001011010001", b"00111010001001111001110101010111"), -- 0.000639399 + 9.93438e-23 = 0.000639399
	(b"10111001101000111111000110100000", b"00000000000000000000000000000000"),
	(b"11010101010011010010000011101100", b"11010101010011010010000011101100"), -- -0.000312698 + -1.40963e+13 = -1.40963e+13
	(b"11010101000101011001111000001111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.02816e+13 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101010010001000000111101010111", b"10101010010001000000111101010111"), -- -0 + -1.74136e-13 = -1.74136e-13
	(b"10011111110010101100000101001100", b"00000000000000000000000000000000"),
	(b"11001011001010010001011110111111", b"11001011001010010001011110111111"), -- -8.58701e-20 + -1.10817e+07 = -1.10817e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011011100001001010001100100000", b"11011011100001001010001100100000"), -- -0 + -7.46681e+16 = -7.46681e+16
	(b"01001100100111001100001100101001", b"00000000000000000000000000000000"),
	(b"01001111110110100100011110010111", b"01001111110111001011101010100100"), -- 8.21886e+07 + 7.32425e+09 = 7.40644e+09
	(b"10101111001111010111100101101000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10101111001111010111100101101000"), -- -1.72326e-10 + -0 = -1.72326e-10
	(b"01110100010100011010010101000010", b"00000000000000000000000000000000"),
	(b"00001100011001000010001101011111", b"01110100010100011010010101000010"), -- 6.64393e+31 + 1.75751e-31 = 6.64393e+31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011001001101110111010100000010", b"11111111100000000000000000000000"), -- -inf + -9.48451e-24 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00010011000111101100111110011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000001010000000", b"00010011000111101100111110011010"), -- 2.00448e-27 + 8.96831e-43 = 2.00448e-27
	(b"01111011000011111111110100010111", b"00000000000000000000000000000000"),
	(b"00110001000011010001000010110100", b"01111011000011111111110100010111"), -- 7.47632e+35 + 2.05277e-09 = 7.47632e+35
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10010010111011101010010100011011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10010010111011101010010100011011"), -- -1.50606e-27 + -0 = -1.50606e-27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10001010101110001001001011100100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10001010101110001001001011100100"), -- -1.77738e-32 + -0 = -1.77738e-32
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11011001011011100110111101010111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.19459e+15 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001100000110000010100001000010", b"10001100000110000010100001000010"), -- -0 + -1.17218e-31 = -1.17218e-31
	(b"01101011101111101000111101101010", b"00000000000000000000000000000000"),
	(b"01011000101011010101101110111100", b"01101011101111101000111101101010"), -- 4.60746e+26 + 1.52488e+15 = 4.60746e+26
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100110001111100110010100000011", b"00100110001111100110010100000011"), -- 0 + 6.60564e-16 = 6.60564e-16
	(b"11111100101011000101001111000000", b"00000000000000000000000000000000"),
	(b"11111011101011000111111011111011", b"11111100110101110111001101111111"), -- -7.15819e+36 + -1.7913e+36 = -8.94949e+36
	(b"11000001100100000001100111000001", b"00000000000000000000000000000000"),
	(b"11010010110111100101001010100101", b"11010010110111100101001010100101"), -- -18.0126 + -4.77435e+11 = -4.77435e+11
	(b"11100111100000100101100100010100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.2311e+24 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000100001100001101000101111101", b"01111111100000000000000000000000"), -- inf + 707.273 = inf
	(b"10010000100101001111101100111111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10010000100101001111101100111111"), -- -5.87628e-29 + -0 = -5.87628e-29
	(b"11101101001110110010100101110000", b"00000000000000000000000000000000"),
	(b"10011111110100000001011110010010", b"11101101001110110010100101110000"), -- -3.62024e+27 + -8.81304e-20 = -3.62024e+27
	(b"11100111010010011111010001000100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -9.53702e+23 + -inf = -inf
	(b"10010001101100100101110010000001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10010001101100100101110010000001"), -- -2.81405e-28 + -0 = -2.81405e-28
	(b"11010000110110101111100011011010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.93899e+10 + -inf = -inf
	(b"01100001001110110001110110111101", b"00000000000000000000000000000000"),
	(b"01011011000001010110101001110100", b"01100001001110110010011000010100"), -- 2.1573e+20 + 3.75532e+16 = 2.15768e+20
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101001101010010010100001000111", b"01111111100000000000000000000000"), -- inf + 7.51209e-14 = inf
	(b"10011001001100011001101100011110", b"00000000000000000000000000000000"),
	(b"11010100111010000110011100001000", b"11010100111010000110011100001000"), -- -9.18201e-24 + -7.98529e+12 = -7.98529e+12
	(b"10111101011011001011101101110011", b"00000000000000000000000000000000"),
	(b"10010001000100001111001111100111", b"10111101011011001011101101110011"), -- -0.057796 + -1.14348e-28 = -0.057796
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111110111100000100111111101111", b"01111110111100000100111111101111"), -- 0 + 1.59715e+38 = 1.59715e+38
	(b"11101100011011000000011011010001", b"00000000000000000000000000000000"),
	(b"11000110100000110101100111010001", b"11101100011011000000011011010001"), -- -1.14135e+27 + -16812.9 = -1.14135e+27
	(b"00111000111100100100100010011010", b"00000000000000000000000000000000"),
	(b"01111001010110011101010110001010", b"01111001010110011101010110001010"), -- 0.00011553 + 7.06912e+34 = 7.06912e+34
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001111101011111110001001001", b"11111111100000000000000000000000"), -- -inf + -3.71723e+25 = -inf
	(b"11000010001001110000011111010111", b"00000000000000000000000000000000"),
	(b"10110101111111001111101000100010", b"11000010001001110000011111010111"), -- -41.7577 + -1.88483e-06 = -41.7577
	(b"10100111010101111001111000110110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100111010101111001111000110110"), -- -2.9923e-15 + -0 = -2.9923e-15
	(b"00000000000000001111111001001111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000001111111001001111"), -- 9.12287e-41 + 0 = 9.12287e-41
	(b"11110010000000000110100001110000", b"00000000000000000000000000000000"),
	(b"11001101110111000000000111110001", b"11110010000000000110100001110000"), -- -2.54338e+30 + -4.61389e+08 = -2.54338e+30
	(b"00010010001010001000111100101111", b"00000000000000000000000000000000"),
	(b"01101111101111111000001011011111", b"01101111101111111000001011011111"), -- 5.31879e-28 + 1.1854e+29 = 1.1854e+29
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110000011010111001110111001101", b"11111111100000000000000000000000"), -- -inf + -2.91679e+29 = -inf
	(b"10000000000000000000000101000001", b"00000000000000000000000000000000"),
	(b"10101011001101101110100001111111", b"10101011001101101110100001111111"), -- -4.49817e-43 + -6.4982e-13 = -6.4982e-13
	(b"10001011111011010101100010010010", b"00000000000000000000000000000000"),
	(b"11101011111111001000111010100110", b"11101011111111001000111010100110"), -- -9.14223e-32 + -6.10646e+26 = -6.10646e+26
	(b"11000110110001111011110110110001", b"00000000000000000000000000000000"),
	(b"10010101001010110000010101100001", b"11000110110001111011110110110001"), -- -25566.8 + -3.45374e-26 = -25566.8
	(b"01010111000110010110001100000110", b"00000000000000000000000000000000"),
	(b"01000011000110011010100110111010", b"01010111000110010110001100000110"), -- 1.68651e+14 + 153.663 = 1.68651e+14
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010100101011101001110010011010", b"11010100101011101001110010011010"), -- -0 + -5.99961e+12 = -5.99961e+12
	(b"10000110100000000001110110011010", b"00000000000000000000000000000000"),
	(b"10110010100001001000011110000011", b"10110010100001001000011110000011"), -- -4.81917e-35 + -1.54284e-08 = -1.54284e-08
	(b"11011110000001100111100110110111", b"00000000000000000000000000000000"),
	(b"10010001100001111101001011000000", b"11011110000001100111100110110111"), -- -2.42249e+18 + -2.14291e-28 = -2.42249e+18
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10101010001011101110111001010100", b"00000000000000000000000000000000"),
	(b"10011001000011111111010010010010", b"10101010001011101110111001010100"), -- -1.5537e-13 + -7.44232e-24 = -1.5537e-13
	(b"00010010100101001111101001110010", b"00000000000000000000000000000000"),
	(b"00000000000000100101001100011101", b"00010010100101001111101001110010"), -- 9.40185e-28 + 2.13486e-40 = 9.40185e-28
	(b"00011111100110101010011001010110", b"00000000000000000000000000000000"),
	(b"01101111001000100110001100101111", b"01101111001000100110001100101111"), -- 6.54967e-20 + 5.02565e+28 = 5.02565e+28
	(b"10011011111101011001001101111111", b"00000000000000000000000000000000"),
	(b"10101111111010111011111001110001", b"10101111111010111011111001110001"), -- -4.06272e-22 + -4.28816e-10 = -4.28816e-10
	(b"11011100010101011101100011101000", b"00000000000000000000000000000000"),
	(b"10110100101000101011111110110110", b"11011100010101011101100011101000"), -- -2.40771e+17 + -3.03143e-07 = -2.40771e+17
	(b"11100000110001111101101001111001", b"00000000000000000000000000000000"),
	(b"11001010000001011001110011100001", b"11100000110001111101101001111001"), -- -1.15208e+20 + -2.18911e+06 = -1.15208e+20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00101101100110111000100011000100", b"00000000000000000000000000000000"),
	(b"01100101100010110100101100010001", b"01100101100010110100101100010001"), -- 1.76822e-11 + 8.22242e+22 = 8.22242e+22
	(b"11001100101101010011100110010110", b"00000000000000000000000000000000"),
	(b"10110110100101101000111001101001", b"11001100101101010011100110010110"), -- -9.50141e+07 + -4.48693e-06 = -9.50141e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00101101110110111001110100001100", b"00000000000000000000000000000000"),
	(b"00001110001000001001111001010011", b"00101101110110111001110100001100"), -- 2.49672e-11 + 1.97978e-30 = 2.49672e-11
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011011001101000000100111000001", b"00011011001101000000100111000001"), -- 0 + 1.48924e-22 = 1.48924e-22
	(b"10000000001001011001001000001110", b"00000000000000000000000000000000"),
	(b"10111010010010100101001010000100", b"10111010010010100101001010000100"), -- -3.45031e-39 + -0.000771798 = -0.000771798
	(b"01100111001111000010011101010111", b"00000000000000000000000000000000"),
	(b"00111010001001111110000011000101", b"01100111001111000010011101010111"), -- 8.88531e+23 + 0.000640404 = 8.88531e+23
	(b"10110010100000101000101101011011", b"00000000000000000000000000000000"),
	(b"10000110011000010111000111010000", b"10110010100000101000101101011011"), -- -1.51974e-08 + -4.24014e-35 = -1.51974e-08
	(b"01100010110110111101010111000010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.02762e+21 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10101101111111101100000111001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10101101111111101100000111001101"), -- -2.89625e-11 + -0 = -2.89625e-11
	(b"11000000011110011110100010001101", b"00000000000000000000000000000000"),
	(b"10011111001110100110011011100011", b"11000000011110011110100010001101"), -- -3.90482 + -3.94721e-20 = -3.90482
	(b"01001011010101101010010111100100", b"00000000000000000000000000000000"),
	(b"01111000000000111100110000011010", b"01111000000000111100110000011010"), -- 1.40672e+07 + 1.06927e+34 = 1.06927e+34
	(b"00010010100111100001000111110111", b"00000000000000000000000000000000"),
	(b"00000011111101110111000000100010", b"00010010100111100001000111110111"), -- 9.97563e-28 + 1.45431e-36 = 9.97563e-28
	(b"00100011110111100000111110100100", b"00000000000000000000000000000000"),
	(b"00011010110011110100011011010010", b"00100011110111100000111111011000"), -- 2.40759e-17 + 8.57276e-23 = 2.4076e-17
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110111000101000110001110010010", b"00110111000101000110001110010010"), -- 0 + 8.84467e-06 = 8.84467e-06
	(b"11011010000001111111010001101011", b"00000000000000000000000000000000"),
	(b"11001000111000101100001101101001", b"11011010000001111111010001101011"), -- -9.56697e+15 + -464411 = -9.56697e+15
	(b"00000101001111111110101000101101", b"00000000000000000000000000000000"),
	(b"01110001011011011011100100010001", b"01110001011011011011100100010001"), -- 9.02379e-36 + 1.17715e+30 = 1.17715e+30
	(b"00100001110000000110001001100100", b"00000000000000000000000000000000"),
	(b"00111011000001101001000100110101", b"00111011000001101001000100110101"), -- 1.30365e-18 + 0.00205333 = 0.00205333
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00110000100010110000101101101100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00110000100010110000101101101100"), -- 1.01168e-09 + 0 = 1.01168e-09
	(b"10110001001101100111000011100010", b"00000000000000000000000000000000"),
	(b"10000101100100101111100011010110", b"10110001001101100111000011100010"), -- -2.65487e-09 + -1.38212e-35 = -2.65487e-09
	(b"01001101100011001010011100010100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.9497e+08 + inf = inf
	(b"01110110000101111011011110010101", b"00000000000000000000000000000000"),
	(b"01010110100011011001010101000000", b"01110110000101111011011110010101"), -- 7.69297e+32 + 7.78361e+13 = 7.69297e+32
	(b"11011111001101010011101111010010", b"00000000000000000000000000000000"),
	(b"10011001010000110111110000101100", b"11011111001101010011101111010010"), -- -1.30593e+19 + -1.01063e-23 = -1.30593e+19
	(b"00110100010000000111110001000010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.79266e-07 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00111111010110111010011110100000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0.858027 + inf = inf
	(b"00001111011000111100100101100001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.12307e-29 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00110011000101111011000010010010", b"00000000000000000000000000000000"),
	(b"00001010001100010010101010001111", b"00110011000101111011000010010010"), -- 3.5318e-08 + 8.53024e-33 = 3.5318e-08
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101001110010010111000000000100", b"11111111100000000000000000000000"), -- -inf + -8.94562e-14 = -inf
	(b"00000111011011001100111011100111", b"00000000000000000000000000000000"),
	(b"00010000000000111000010101011111", b"00010000000000111000010110011010"), -- 1.78155e-34 + 2.59379e-29 = 2.59381e-29
	(b"11001010100101001001011000010111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001010100101001001011000010111"), -- -4.86888e+06 + -0 = -4.86888e+06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11000000100110010110111010011001", b"00000000000000000000000000000000"),
	(b"11010010100101100100010000010111", b"11010010100101100100010000010111"), -- -4.79475 + -3.22694e+11 = -3.22694e+11
	(b"01100100000110010111001111011000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.13228e+22 + inf = inf
	(b"10111110000000110001010010101011", b"00000000000000000000000000000000"),
	(b"11101000010111011110001011101011", b"11101000010111011110001011101011"), -- -0.128009 + -4.19132e+24 = -4.19132e+24
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111001001001111001011101010001", b"11111111100000000000000000000000"), -- -inf + -5.43864e+34 = -inf
	(b"10011010011001100100101101111100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10011010011001100100101101111100"), -- -4.76239e-23 + -0 = -4.76239e-23
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001010011110101001100111101001", b"01111111100000000000000000000000"), -- inf + 4.10585e+06 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111010110001001101101010111110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.11063e+35 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011111110110111111000111110001", b"11111111100000000000000000000000"), -- -inf + -3.16974e+19 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110111101100111000101011000011", b"11111111100000000000000000000000"), -- -inf + -7.28309e+33 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111010111110101010011111010111", b"11111111100000000000000000000000"), -- -inf + -6.50739e+35 = -inf
	(b"00111000001001101110111010111100", b"00000000000000000000000000000000"),
	(b"01101110101101000100101111010000", b"01101110101101000100101111010000"), -- 3.97998e-05 + 2.78995e+28 = 2.78995e+28
	(b"00111100101000100001000101101001", b"00000000000000000000000000000000"),
	(b"01011100100010101111001000001011", b"01011100100010101111001000001011"), -- 0.0197837 + 3.12877e+17 = 3.12877e+17
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101110101100101000000100111011", b"00101110101100101000000100111011"), -- 0 + 8.11746e-11 = 8.11746e-11
	(b"01011000010111000011011110110101", b"00000000000000000000000000000000"),
	(b"01100010101110110001001001100011", b"01100010101110110001001001101010"), -- 9.68527e+14 + 1.72543e+21 = 1.72543e+21
	(b"00010110010111010111000110010100", b"00000000000000000000000000000000"),
	(b"01100100000111011100101110100001", b"01100100000111011100101110100001"), -- 1.78881e-25 + 1.16432e+22 = 1.16432e+22
	(b"11000101100111000111010110001011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000101100111000111010110001011"), -- -5006.69 + -0 = -5006.69
	(b"00001001110110101110110100111100", b"00000000000000000000000000000000"),
	(b"01011001001100010011100100111101", b"01011001001100010011100100111101"), -- 5.27047e-33 + 3.11775e+15 = 3.11775e+15
	(b"11110000001100110100101010010001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.21952e+29 + -inf = -inf
	(b"00000111110001111001011010111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000111011010", b"00000111110001111001011010111011"), -- 3.00308e-34 + 6.64215e-43 = 3.00308e-34
	(b"10000000000000001001000110000100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.22012e-41 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001110100100001001000000010101", b"10001110100100001001000000010101"), -- -0 + -3.56375e-30 = -3.56375e-30
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100100110100111111111010000111", b"11111111100000000000000000000000"), -- -inf + -9.19378e-17 = -inf
	(b"11011110101000010011010000001001", b"00000000000000000000000000000000"),
	(b"11111001100011101001010011001101", b"11111001100011101001010011001101"), -- -5.80796e+18 + -9.25405e+34 = -9.25405e+34
	(b"00110010000000011010000011100101", b"00000000000000000000000000000000"),
	(b"00111111000010101100011111010100", b"00111111000010101100011111010100"), -- 7.54537e-09 + 0.542112 = 0.542112
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11101010010010111010010000100110", b"00000000000000000000000000000000"),
	(b"10110100010011011110111110100110", b"11101010010010111010010000100110"), -- -6.15468e+25 + -1.91793e-07 = -6.15468e+25
	(b"10010101110100010100101000101111", b"00000000000000000000000000000000"),
	(b"11101000101111110001010111010001", b"11101000101111110001010111010001"), -- -8.45315e-26 + -7.219e+24 = -7.219e+24
	(b"10111110010001111001110001001111", b"00000000000000000000000000000000"),
	(b"11011010100000111000101000000101", b"11011010100000111000101000000101"), -- -0.194932 + -1.85125e+16 = -1.85125e+16
	(b"10110001100101000000100001001100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110001100101000000100001001100"), -- -4.30831e-09 + -0 = -4.30831e-09
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101110100100001100100001010011", b"01101110100100001100100001010011"), -- 0 + 2.2404e+28 = 2.2404e+28
	(b"10000001110011110111110110100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000001110011110111110110100110"), -- -7.62201e-38 + -0 = -7.62201e-38
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000010110111010", b"11111111100000000000000000000000"), -- -inf + -2.0543e-42 = -inf
	(b"01000010001010100111100011000111", b"00000000000000000000000000000000"),
	(b"01011001001101010000101100010110", b"01011001001101010000101100010110"), -- 42.6179 + 3.18495e+15 = 3.18495e+15
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001111011010011110100101110000", b"01111111100000000000000000000000"), -- inf + 1.15327e-29 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001001000110111101011101101110", b"11111111100000000000000000000000"), -- -inf + -638327 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101100101111011000101010110011", b"01111111100000000000000000000000"), -- inf + 1.83314e+27 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01101001000011011000011000010000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101001000011011000011000010000"), -- 1.06932e+25 + 0 = 1.06932e+25
	(b"11011010111101110011111110001011", b"00000000000000000000000000000000"),
	(b"10000000001111011010000010100100", b"11011010111101110011111110001011"), -- -3.47971e+16 + -5.65959e-39 = -3.47971e+16
	(b"00111001100110111110001110010110", b"00000000000000000000000000000000"),
	(b"00011110001011010001101000111100", b"00111001100110111110001110010110"), -- 0.000297335 + 9.16397e-21 = 0.000297335
	(b"00101110001010001000001000000101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00101110001010001000001000000101"), -- 3.83143e-11 + 0 = 3.83143e-11
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011001100100100100100101101110", b"10011001100100100100100101101110"), -- -0 + -1.51257e-23 = -1.51257e-23
	(b"00100100010111101100001000011000", b"00000000000000000000000000000000"),
	(b"00010010110111101001000011111010", b"00100100010111101100001000011000"), -- 4.8303e-17 + 1.40459e-27 = 4.8303e-17
	(b"11011110110101011000110000100010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11011110110101011000110000100010"), -- -7.69386e+18 + -0 = -7.69386e+18
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100000011010111001101111110101", b"11111111100000000000000000000000"), -- -inf + -6.79097e+19 = -inf
	(b"11111101100000110001101111110101", b"00000000000000000000000000000000"),
	(b"11000110100000001101111101100010", b"11111101100000110001101111110101"), -- -2.17843e+37 + -16495.7 = -2.17843e+37
	(b"11110100000101100111001110000001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.76799e+31 + -inf = -inf
	(b"01000101110010101010000100001011", b"00000000000000000000000000000000"),
	(b"00111101100111011101111111100010", b"01000101110010101010000110101001"), -- 6484.13 + 0.0770872 = 6484.21
	(b"10011000011001100110100110111101", b"00000000000000000000000000000000"),
	(b"11010111001010011010000100110000", b"11010111001010011010000100110000"), -- -2.97802e-24 + -1.8651e+14 = -1.8651e+14
	(b"00111101100001010000011010111111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111101100001010000011010111111"), -- 0.0649543 + 0 = 0.0649543
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010001100010100100101010110001", b"11010001100010100100101010110001"), -- -0 + -7.42448e+10 = -7.42448e+10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11011011100101110110011000000010", b"00000000000000000000000000000000"),
	(b"10011010111110011000000100001100", b"11011011100101110110011000000010"), -- -8.52298e+16 + -1.03192e-22 = -8.52298e+16
	(b"10000000000000000000011010111101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000011010111101"), -- -2.41724e-42 + -0 = -2.41724e-42
	(b"10000000000000000000000000010010", b"00000000000000000000000000000000"),
	(b"11000101000010101110100000100111", b"11000101000010101110100000100111"), -- -2.52234e-44 + -2222.51 = -2222.51
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111010011110010010111010110001", b"11111111100000000000000000000000"), -- -inf + -0.000950555 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110010011110011111011011110100", b"11110010011110011111011011110100"), -- -0 + -4.95106e+30 = -4.95106e+30
	(b"10000101010110011101001011000000", b"00000000000000000000000000000000"),
	(b"10100111000000000100111001000011", b"10100111000000000100111001000011"), -- -1.0242e-35 + -1.7806e-15 = -1.7806e-15
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101110111000111011001101010111", b"01111111100000000000000000000000"), -- inf + 1.03546e-10 = inf
	(b"00110010110001011100011101011011", b"00000000000000000000000000000000"),
	(b"00100001101110001011110100001100", b"00110010110001011100011101011011"), -- 2.30245e-08 + 1.25184e-18 = 2.30245e-08
	(b"10101001010001100011010010000110", b"00000000000000000000000000000000"),
	(b"10000010001000100101010111001111", b"10101001010001100011010010000110"), -- -4.40104e-14 + -1.19265e-37 = -4.40104e-14
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000111011101101110100", b"10000000000000111011101101110100"), -- -0 + -3.42752e-40 = -3.42752e-40
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101011011110001000101000100100", b"11101011011110001000101000100100"), -- -0 + -3.00466e+26 = -3.00466e+26
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000011100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000011100"), -- 3.92364e-44 + 0 = 3.92364e-44
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000001000001010010100000011", b"00000000000000000000000000000000"),
	(b"00110101001000011111000011000010", b"00110101001000011111000011000010"), -- 2.99793e-39 + 6.03275e-07 = 6.03275e-07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000111010011010011", b"00000000000000000111010011010011"), -- 0 + 4.19086e-41 = 4.19086e-41
	(b"10010110010101011110000101011001", b"00000000000000000000000000000000"),
	(b"11000010111001100101000000001100", b"11000010111001100101000000001100"), -- -1.72771e-25 + -115.156 = -115.156
	(b"01101010100001111000000010000110", b"00000000000000000000000000000000"),
	(b"01111001110000000110010100001010", b"01111001110000000110010100001010"), -- 8.1906e+25 + 1.24871e+35 = 1.24871e+35
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11000100100010010000110010001000", b"00000000000000000000000000000000"),
	(b"11111010001101010001111011000100", b"11111010001101010001111011000100"), -- -1096.39 + -2.35107e+35 = -2.35107e+35
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000101100111111", b"01111111100000000000000000000000"), -- inf + 4.03434e-42 = inf
	(b"01110011101000110001111011010101", b"00000000000000000000000000000000"),
	(b"01011011101001000111001110101101", b"01110011101000110001111011010101"), -- 2.58475e+31 + 9.25782e+16 = 2.58475e+31
	(b"00101000111011010110110111110111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00101000111011010110110111110111"), -- 2.636e-14 + 0 = 2.636e-14
	(b"00011001000100001101111000011101", b"00000000000000000000000000000000"),
	(b"01000101101101101011001101010011", b"01000101101101101011001101010011"), -- 7.48948e-24 + 5846.42 = 5846.42
	(b"00000000000000100100000101111101", b"00000000000000000000000000000000"),
	(b"01000001100110011111011010011011", b"01000001100110011111011010011011"), -- 2.07164e-40 + 19.2454 = 19.2454
	(b"01001011100010110000101000001000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.82241e+07 + inf = inf
	(b"00000000000010001011011110000000", b"00000000000000000000000000000000"),
	(b"01110111101110001111101000101011", b"01110111101110001111101000101011"), -- 8.00511e-40 + 7.50357e+33 = 7.50357e+33
	(b"11100110010101000010001110010110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11100110010101000010001110010110"), -- -2.5045e+23 + -0 = -2.5045e+23
	(b"10111100010000000001011000100001", b"00000000000000000000000000000000"),
	(b"11100111100000010101010001100011", b"11100111100000010101010001100011"), -- -0.011724 + -1.22148e+24 = -1.22148e+24
	(b"11100100111011000100100001110100", b"00000000000000000000000000000000"),
	(b"10011110110001011101110111000011", b"11100100111011000100100001110100"), -- -3.48692e+22 + -2.09499e-20 = -3.48692e+22
	(b"01011001010000101010110101001011", b"00000000000000000000000000000000"),
	(b"00110100110101100001001011011010", b"01011001010000101010110101001011"), -- 3.42479e+15 + 3.98743e-07 = 3.42479e+15
	(b"11010100011010010100000001000001", b"00000000000000000000000000000000"),
	(b"11011000000011001001100011110100", b"11011000000011011000001000110100"), -- -4.00722e+12 + -6.18354e+14 = -6.22361e+14
	(b"10101110011111011000101110110111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10101110011111011000101110110111"), -- -5.76496e-11 + -0 = -5.76496e-11
	(b"01010101110110111001011111001101", b"00000000000000000000000000000000"),
	(b"00000000000000000111111100010100", b"01010101110110111001011111001101"), -- 3.01806e+13 + 4.5587e-41 = 3.01806e+13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000111100011101111100110000000", b"11111111100000000000000000000000"), -- -inf + -73203 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001110101010000010001001000", b"11101001110101010000010001001000"), -- -0 + -3.21902e+25 = -3.21902e+25
	(b"01110110111101110101001110011000", b"00000000000000000000000000000000"),
	(b"00111101010010011000000000000001", b"01110110111101110101001110011000"), -- 2.50819e+33 + 0.0491943 = 2.50819e+33
	(b"11100101101011110111111100111111", b"00000000000000000000000000000000"),
	(b"10010111100011000111111100001110", b"11100101101011110111111100111111"), -- -1.03595e+23 + -9.07936e-25 = -1.03595e+23
	(b"11111001110100000000000100100011", b"00000000000000000000000000000000"),
	(b"10110101001101001100011110100011", b"11111001110100000000000100100011"), -- -1.35003e+35 + -6.73457e-07 = -1.35003e+35
	(b"10111101010101000111011011011000", b"00000000000000000000000000000000"),
	(b"11110000100011110100001110100110", b"11110000100011110100001110100110"), -- -0.0518712 + -3.54705e+29 = -3.54705e+29
	(b"00100011000111100101111111110001", b"00000000000000000000000000000000"),
	(b"01010110000000000000001000010101", b"01010110000000000000001000010101"), -- 8.58551e-18 + 3.51866e+13 = 3.51866e+13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10100000100000100011100011001000", b"00000000000000000000000000000000"),
	(b"11011001111011011010001010110001", b"11011001111011011010001010110001"), -- -2.20604e-19 + -8.36106e+15 = -8.36106e+15
	(b"00011101011100011010000011101100", b"00000000000000000000000000000000"),
	(b"01111101001010001110101101000110", b"01111101001010001110101101000110"), -- 3.19793e-21 + 1.40332e+37 = 1.40332e+37
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000010010111", b"11111111100000000000000000000000"), -- -inf + -2.11596e-43 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011101101101101101101010010101", b"11111111100000000000000000000000"), -- -inf + -4.8401e-21 = -inf
	(b"00101111010000111111010011100001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.78221e-10 + inf = inf
	(b"10111100101010110001001111011000", b"00000000000000000000000000000000"),
	(b"10101000011010110100101111010000", b"10111100101010110001001111011000"), -- -0.0208835 + -1.30616e-14 = -0.0208835
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011100000100101110000011100110", b"01111111100000000000000000000000"), -- inf + 4.8598e-22 = inf
	(b"00000100111000101111101001100101", b"00000000000000000000000000000000"),
	(b"01010100001100001111110101000100", b"01010100001100001111110101000100"), -- 5.33623e-36 + 3.04065e+12 = 3.04065e+12
	(b"11000001111010010101101110001101", b"00000000000000000000000000000000"),
	(b"11011110001101010111110000111111", b"11011110001101010111110000111111"), -- -29.1697 + -3.26935e+18 = -3.26935e+18
	(b"10110111010100011001110011011010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.24939e-05 + -inf = -inf
	(b"10000000000000000000000000010100", b"00000000000000000000000000000000"),
	(b"11111101111001001111110011111111", b"11111101111001001111110011111111"), -- -2.8026e-44 + -3.80472e+37 = -3.80472e+37
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01011011111100110111101100101101", b"00000000000000000000000000000000"),
	(b"00111011010000010011110011101000", b"01011011111100110111101100101101"), -- 1.37068e+17 + 0.00294858 = 1.37068e+17
	(b"10111010101111111001100011001100", b"00000000000000000000000000000000"),
	(b"11010111101110111010000100100100", b"11010111101110111010000100100100"), -- -0.00146177 + -4.12602e+14 = -4.12602e+14
	(b"00110111011000111101110010100010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.35816e-05 + inf = inf
	(b"01100000100110110011100010110001", b"00000000000000000000000000000000"),
	(b"01001100001010011110010101011101", b"01100000100110110011100010110001"), -- 8.94791e+19 + 4.45372e+07 = 8.94791e+19
	(b"10000000000000000000101001110100", b"00000000000000000000000000000000"),
	(b"11000100111011110110111111101010", b"11000100111011110110111111101010"), -- -3.74987e-42 + -1915.5 = -1915.5
	(b"00110001010110000110101110010100", b"00000000000000000000000000000000"),
	(b"01010111001010011010111110011010", b"01010111001010011010111110011010"), -- 3.14933e-09 + 1.86572e+14 = 1.86572e+14
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00101111110101100100010100100111", b"00000000000000000000000000000000"),
	(b"01101010000011110100010010011100", b"01101010000011110100010010011100"), -- 3.89755e-10 + 4.33001e+25 = 4.33001e+25
	(b"11011001011100111000101000100001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.28439e+15 + -inf = -inf
	(b"10000000000000000000000111011111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.71222e-43 + -inf = -inf
	(b"10010010100011111110100101110011", b"00000000000000000000000000000000"),
	(b"11000111100100000101011001001010", b"11000111100100000101011001001010"), -- -9.08212e-28 + -73900.6 = -73900.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000101110100110101110101010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.98766e-35 + -inf = -inf
	(b"10100111000001000100011000101010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.83567e-15 + -inf = -inf
	(b"00111001011010000011000101100111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111001011010000011000101100111"), -- 0.000221436 + 0 = 0.000221436
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10010011100001010101010001100011", b"00000000000000000000000000000000"),
	(b"10100111100000110011001010101111", b"10100111100000110011001010101111"), -- -3.36571e-27 + -3.64148e-15 = -3.64148e-15
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010101111110011011100100110000", b"01111111100000000000000000000000"), -- inf + 3.43217e+13 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000111111", b"10000000000000000000000000111111"), -- -0 + -8.82818e-44 = -8.82818e-44
	(b"01101000001100000110100001110000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101000001100000110100001110000"), -- 3.33225e+24 + 0 = 3.33225e+24
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001011100010010100100100100011", b"10001011100010010100100100100011"), -- -0 + -5.28805e-32 = -5.28805e-32
	(b"10101011100001000011010101110101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -9.394e-13 + -inf = -inf
	(b"10110000000110001001110111100110", b"00000000000000000000000000000000"),
	(b"11110110101000011011000110110010", b"11110110101000011011000110110010"), -- -5.55217e-10 + -1.63977e+33 = -1.63977e+33
	(b"11011010110001010110001111001101", b"00000000000000000000000000000000"),
	(b"10101100101100101100101110100100", b"11011010110001010110001111001101"), -- -2.77802e+16 + -5.08167e-12 = -2.77802e+16
	(b"01111001111110101110101010100100", b"00000000000000000000000000000000"),
	(b"00101101011101000001001011001000", b"01111001111110101110101010100100"), -- 1.62854e+35 + 1.3874e-11 = 1.62854e+35
	(b"00010100110001000111110001010100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.984e-26 + inf = inf
	(b"01010011101111011100101101001010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.63032e+12 + inf = inf
	(b"01100110001011011011100101000100", b"00000000000000000000000000000000"),
	(b"01010111110001100010110011101010", b"01100110001011011011100101000100"), -- 2.05097e+23 + 4.35792e+14 = 2.05097e+23
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11000000101101010010110010000000", b"00000000000000000000000000000000"),
	(b"10000100101111110101100111000110", b"11000000101101010010110010000000"), -- -5.66168 + -4.49863e-36 = -5.66168
	(b"00100111100011011100010001010010", b"00000000000000000000000000000000"),
	(b"01000011101111001110101001000100", b"01000011101111001110101001000100"), -- 3.93482e-15 + 377.83 = 377.83
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01010110100000110111111100111011", b"00000000000000000000000000000000"),
	(b"00010010000111111000001011101110", b"01010110100000110111111100111011"), -- 7.22912e+13 + 5.03329e-28 = 7.22912e+13
	(b"01111010110101110000000100111101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.58184e+35 + inf = inf
	(b"00110000110110100110101101110110", b"00000000000000000000000000000000"),
	(b"01101101000000110100001111111010", b"01101101000000110100001111111010"), -- 1.58921e-09 + 2.53904e+27 = 2.53904e+27
	(b"11110101110010111011000011110101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.16419e+32 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011000011110111111111000101111", b"01011000011110111111111000101111"), -- 0 + 1.10828e+15 = 1.10828e+15
	(b"00000100011011101010011100101011", b"00000000000000000000000000000000"),
	(b"01000010001110010011111100001011", b"01000010001110010011111100001011"), -- 2.80535e-36 + 46.3116 = 46.3116
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000101011011101110001000101101", b"11111111100000000000000000000000"), -- -inf + -3822.14 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110001001110000110", b"00111111101100110001001110000110"), -- 0 + 1.39903 = 1.39903
	(b"01111000001001110010101100111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111000001001110010101100111011"), -- 1.35623e+34 + 0 = 1.35623e+34
	(b"11111000100110111010011100110100", b"00000000000000000000000000000000"),
	(b"10011111001000010100001101100101", b"11111000100110111010011100110100"), -- -2.52562e+34 + -3.41488e-20 = -2.52562e+34
	(b"10000000000000000000000000100010", b"00000000000000000000000000000000"),
	(b"11111111000110011100110010100000", b"11111111000110011100110010100000"), -- -4.76441e-44 + -2.04434e+38 = -2.04434e+38
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011110100101011000110001011100", b"00011110100101011000110001011100"), -- 0 + 1.5834e-20 = 1.5834e-20
	(b"00000000001100110001001110011010", b"00000000000000000000000000000000"),
	(b"01100101101010001001101001110100", b"01100101101010001001101001110100"), -- 4.69064e-39 + 9.95258e+22 = 9.95258e+22
	(b"11100000110000101110010011101001", b"00000000000000000000000000000000"),
	(b"11111011100111111110000011111000", b"11111011100111111110000011111000"), -- -1.12349e+20 + -1.66028e+36 = -1.66028e+36
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01001011101000001110010101011011", b"00000000000000000000000000000000"),
	(b"01001000111110000110101001110000", b"01001011101001001100011100000101"), -- 2.1089e+07 + 508756 = 2.15977e+07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000001110111001100111001101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000001110111001100111001101"), -- 5.47347e-39 + 0 = 5.47347e-39
	(b"10101000110001000110110001101000", b"00000000000000000000000000000000"),
	(b"10111100100100100000100000110101", b"10111100100100100000100000110101"), -- -2.18074e-14 + -0.0178262 = -0.0178262
	(b"11000100101010100001011001000001", b"00000000000000000000000000000000"),
	(b"11110010001001001001001000111001", b"11110010001001001001001000111001"), -- -1360.7 + -3.25967e+30 = -3.25967e+30
	(b"00001101101011110100010100101011", b"00000000000000000000000000000000"),
	(b"00110001110110010111101001000010", b"00110001110110010111101001000010"), -- 1.08019e-30 + 6.32943e-09 = 6.32943e-09
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01000110101011000010000101010100", b"00000000000000000000000000000000"),
	(b"01011111100111010010110001011100", b"01011111100111010010110001011100"), -- 22032.7 + 2.26511e+19 = 2.26511e+19
	(b"00010110100000011100001010101001", b"00000000000000000000000000000000"),
	(b"00010101110010010101001011001110", b"00010110101101000001011101011100"), -- 2.09639e-25 + 8.13139e-26 = 2.90953e-25
	(b"01100111100101101011011110100101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.42349e+24 + inf = inf
	(b"10110101101101100010110000100100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.35729e-06 + -inf = -inf
	(b"11111100111000010010110011111111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -9.35344e+36 + -inf = -inf
	(b"10110100111111000101010111111110", b"00000000000000000000000000000000"),
	(b"11011001011010110011000000110011", b"11011001011010110011000000110011"), -- -4.70012e-07 + -4.13748e+15 = -4.13748e+15
	(b"11100001011011010111111011010010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.73814e+20 + -inf = -inf
	(b"10110110101000010000000001001110", b"00000000000000000000000000000000"),
	(b"10101000100000010101011000111110", b"10110110101000010000000001001110"), -- -4.79821e-06 + -1.43593e-14 = -4.79821e-06
	(b"01001101110110010000100001110001", b"00000000000000000000000000000000"),
	(b"00011110101000000110010110101111", b"01001101110110010000100001110001"), -- 4.55151e+08 + 1.69827e-20 = 4.55151e+08
	(b"00001100110001100000110111001100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00001100110001100000110111001100"), -- 3.0515e-31 + 0 = 3.0515e-31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010110000110000101001101001100", b"11111111100000000000000000000000"), -- -inf + -1.23047e-25 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01101010100100100011101100001101", b"00000000000000000000000000000000"),
	(b"00100010100010011101000110010101", b"01101010100100100011101100001101"), -- 8.8391e+25 + 3.73558e-18 = 8.8391e+25
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011000101011110010111111101000", b"00011000101011110010111111101000"), -- 0 + 4.52848e-24 = 4.52848e-24
	(b"00001100100001010001001000010100", b"00000000000000000000000000000000"),
	(b"00010111001100011011110101100010", b"00010111001100011011110101100110"), -- 2.05028e-31 + 5.74308e-25 = 5.74308e-25
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011011100000101011111100001110", b"10011011100000101011111100001110"), -- -0 + -2.16302e-22 = -2.16302e-22
	(b"10100110101000010101100010010000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100110101000010101100010010000"), -- -1.11956e-15 + -0 = -1.11956e-15
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110001011011011001101011100101", b"01111111100000000000000000000000"), -- inf + 1.17656e+30 = inf
	(b"11000010011110010101100000100011", b"00000000000000000000000000000000"),
	(b"10000000111111111111100010110100", b"11000010011110010101100000100011"), -- -62.3361 + -2.35073e-38 = -62.3361
	(b"10101001010101010000111100101010", b"00000000000000000000000000000000"),
	(b"11100110100010011110111111000001", b"11100110100010011110111111000001"), -- -4.73087e-14 + -3.25693e+23 = -3.25693e+23
	(b"10101000011011111111010101011101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.33204e-14 + -inf = -inf
	(b"00000000000000000000000100110011", b"00000000000000000000000000000000"),
	(b"00000000000001100100001000111100", b"00000000000001100100001101101111"), -- 4.30199e-43 + 5.74773e-40 = 5.75204e-40
	(b"11111101111111000000101000111000", b"00000000000000000000000000000000"),
	(b"10000111100100101111010010011011", b"11111101111111000000101000111000"), -- -4.18773e+37 + -2.21114e-34 = -4.18773e+37
	(b"11100000110111011101011001000101", b"00000000000000000000000000000000"),
	(b"10000000000000000011010101100000", b"11100000110111011101011001000101"), -- -1.2788e+20 + -1.91473e-41 = -1.2788e+20
	(b"11010100100010000000001000001011", b"00000000000000000000000000000000"),
	(b"11000110011100101001110001010100", b"11010100100010000000001000001011"), -- -4.6732e+12 + -15527.1 = -4.6732e+12
	(b"01110010000010101011101110101001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01110010000010101011101110101001"), -- 2.74789e+30 + 0 = 2.74789e+30
	(b"00000000000000000000000001111000", b"00000000000000000000000000000000"),
	(b"01010110001110001010000110010011", b"01010110001110001010000110010011"), -- 1.68156e-43 + 5.0751e+13 = 5.0751e+13
	(b"10001110110011001011010001101011", b"00000000000000000000000000000000"),
	(b"11010001111111011011001101010010", b"11010001111111011011001101010010"), -- -5.04636e-30 + -1.36204e+11 = -1.36204e+11
	(b"00101001100100101000110010100011", b"00000000000000000000000000000000"),
	(b"01101101010100100111011011110011", b"01101101010100100111011011110011"), -- 6.5081e-14 + 4.07098e+27 = 4.07098e+27
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101111000000000101111110111111", b"11111111100000000000000000000000"), -- -inf + -1.16755e-10 = -inf
	(b"01001111110000101011110000111110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.53423e+09 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110100001101101100111011101010", b"10110100001101101100111011101010"), -- -0 + -1.70253e-07 = -1.70253e-07
	(b"00111001011110101101110010000001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0.00023924 + inf = inf
	(b"11101000110100100110100011011001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.94905e+24 + -inf = -inf
	(b"10111000111101011111111111100000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0.000117302 + -inf = -inf
	(b"10100101101110000101110111100011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.19825e-16 + -inf = -inf
	(b"10110011001101111000001111111010", b"00000000000000000000000000000000"),
	(b"11110101101100111100101100111110", b"11110101101100111100101100111110"), -- -4.2728e-08 + -4.55832e+32 = -4.55832e+32
	(b"10110110100101001111110000100000", b"00000000000000000000000000000000"),
	(b"10011111000000100101110000101100", b"10110110100101001111110000100000"), -- -4.44009e-06 + -2.76048e-20 = -4.44009e-06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010011100010000001010111111111", b"10010011100010000001010111111111"), -- -0 + -3.43529e-27 = -3.43529e-27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000110010101000010101010101101", b"11000110010101000010101010101101"), -- -0 + -13578.7 = -13578.7
	(b"10001011111011011010010000101110", b"00000000000000000000000000000000"),
	(b"11000001101000000100110100001100", b"11000001101000000100110100001100"), -- -9.15361e-32 + -20.0376 = -20.0376
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111101111001010101001000001000", b"00000000000000000000000000000000"),
	(b"10111111011010011100010011101000", b"11111101111001010101001000001000"), -- -3.81024e+37 + -0.913161 = -3.81024e+37
	(b"01001101111010101010000010000001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.92048e+08 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001101001101111001100011000110", b"11111111100000000000000000000000"), -- -inf + -1.92515e+08 = -inf
	(b"00000010110100000010101000000010", b"00000000000000000000000000000000"),
	(b"01111101100010101110011111000101", b"01111101100010101110011111000101"), -- 3.0587e-37 + 2.30796e+37 = 2.30796e+37
	(b"01001000111011110110110001001011", b"00000000000000000000000000000000"),
	(b"01100011100010001100011011110001", b"01100011100010001100011011110001"), -- 490338 + 5.04618e+21 = 5.04618e+21
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011001000010011111001101100110", b"10011001000010011111001101100110"), -- -0 + -7.13189e-24 = -7.13189e-24
	(b"11010011010001011101001101000100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.49653e+11 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110110010101101011101111011100", b"11111111100000000000000000000000"), -- -inf + -1.08883e+33 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100011110010110010010001", b"11000000100011110010110010010001"), -- -0 + -4.47419 = -4.47419
	(b"01110010111100010011110010110101", b"00000000000000000000000000000000"),
	(b"00110001011101110101101111110001", b"01110010111100010011110010110101"), -- 9.55639e+30 + 3.59955e-09 = 9.55639e+30
	(b"01101100011110000000111110000010", b"00000000000000000000000000000000"),
	(b"00100111011101100110010111001001", b"01101100011110000000111110000010"), -- 1.19955e+27 + 3.41945e-15 = 1.19955e+27
	(b"01101110101101111110010000110110", b"00000000000000000000000000000000"),
	(b"01100100111101110011111010110011", b"01101110101101111110010001000101"), -- 2.84558e+28 + 3.64869e+22 = 2.84559e+28
	(b"00110001100001000110000000010111", b"00000000000000000000000000000000"),
	(b"01001010001110011111000001111111", b"01001010001110011111000001111111"), -- 3.85263e-09 + 3.04643e+06 = 3.04643e+06
	(b"10000010011100100001011011010101", b"00000000000000000000000000000000"),
	(b"11111000000011110011001000010100", b"11111000000011110011001000010100"), -- -1.77859e-37 + -1.16174e+34 = -1.16174e+34
	(b"01010000000111101101001010000101", b"00000000000000000000000000000000"),
	(b"01010010100011000011011111000001", b"01010010100100010010111001010101"), -- 1.06584e+10 + 3.01115e+11 = 3.11774e+11
	(b"11100000010101001111101001010011", b"00000000000000000000000000000000"),
	(b"10101110101100111001000110001011", b"11100000010101001111101001010011"), -- -6.13867e+19 + -8.16583e-11 = -6.13867e+19
	(b"10000000101110001110101011010111", b"00000000000000000000000000000000"),
	(b"11101110110100010001111111110110", b"11101110110100010001111111110110"), -- -1.6982e-38 + -3.23605e+28 = -3.23605e+28
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001000001001000101011101101111", b"11001000001001000101011101101111"), -- -0 + -168286 = -168286
	(b"01101101101110011101001010011110", b"00000000000000000000000000000000"),
	(b"00001000101101000011111000100111", b"01101101101110011101001010011110"), -- 7.18867e+27 + 1.0848e-33 = 7.18867e+27
	(b"10110011000011110010100101011101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000001", b"10110011000011110010100101011101"), -- -3.33324e-08 + -1.4013e-45 = -3.33324e-08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001010111110100011011", b"01111111100000000000000000000000"), -- inf + 5.04057e-40 = inf
	(b"10000000010010100010010101100101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.80924e-39 + -inf = -inf
	(b"11101111000001100111001000000000", b"00000000000000000000000000000000"),
	(b"11001000110111000001111111011110", b"11101111000001100111001000000000"), -- -4.16088e+28 + -450815 = -4.16088e+28
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110010101110010110110100100011", b"10110010101110010110110100100011"), -- -0 + -2.15865e-08 = -2.15865e-08
	(b"10000000111001000011001000110111", b"00000000000000000000000000000000"),
	(b"10101111110011010000110111101001", b"10101111110011010000110111101001"), -- -2.09565e-38 + -3.72992e-10 = -3.72992e-10
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000111100001001100010111100011", b"01111111100000000000000000000000"), -- inf + 67979.8 = inf
	(b"10000011101101101010110001110001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.07366e-36 + -inf = -inf
	(b"00000000000001001001100110110100", b"00000000000000000000000000000000"),
	(b"01101110101100101101111101100011", b"01101110101100101101111101100011"), -- 4.2248e-40 + 2.76792e+28 = 2.76792e+28
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011001100110110111101100000111", b"01011001100110110111101100000111"), -- 0 + 5.47049e+15 = 5.47049e+15
	(b"10000111010010111110101110011111", b"00000000000000000000000000000000"),
	(b"11000110011101001100111110011100", b"11000110011101001100111110011100"), -- -1.53413e-34 + -15667.9 = -15667.9
	(b"01110001011100101001110010000101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.20135e+30 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100101011010111110001001110011", b"10100101011010111110001001110011"), -- -0 + -2.04597e-16 = -2.04597e-16
	(b"11010010100101001000111000100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11010010100101001000111000100110"), -- -3.1902e+11 + -0 = -3.1902e+11
	(b"10000011101100000111101101000100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.03727e-36 + -inf = -inf
	(b"00101111001001011000011001110000", b"00000000000000000000000000000000"),
	(b"01110001101011010010111011000110", b"01110001101011010010111011000110"), -- 1.50544e-10 + 1.71512e+30 = 1.71512e+30
	(b"01011110110101001011000011000101", b"00000000000000000000000000000000"),
	(b"01101010000010000110110010100110", b"01101010000010000110110010101000"), -- 7.66298e+18 + 4.12317e+25 = 4.12318e+25
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001110000010001011011000110010", b"01111111100000000000000000000000"), -- inf + 5.7341e+08 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010000100000000010011011101100", b"11111111100000000000000000000000"), -- -inf + -5.05471e-29 = -inf
	(b"01110010000100100100110101100100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.89782e+30 + inf = inf
	(b"11000010010000111101001101110100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -48.9565 + -inf = -inf
	(b"01101111111010111011001010011001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101111111010111011001010011001"), -- 1.4589e+29 + 0 = 1.4589e+29
	(b"01000100111110000001011101011111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1984.73 + inf = inf
	(b"11110100110100011000100011101111", b"00000000000000000000000000000000"),
	(b"10101110001100110101101000001110", b"11110100110100011000100011101111"), -- -1.32809e+32 + -4.07799e-11 = -1.32809e+32
	(b"01100011000110110001011110101110", b"00000000000000000000000000000000"),
	(b"01010111010101110011011111111011", b"01100011000110110001011110101111"), -- 2.86095e+21 + 2.36635e+14 = 2.86095e+21
	(b"00000000000000111001000001111001", b"00000000000000000000000000000000"),
	(b"00111110010111101010100000110001", b"00111110010111101010100000110001"), -- 3.27334e-40 + 0.217438 = 0.217438
	(b"11011110101110101010001101110001", b"00000000000000000000000000000000"),
	(b"10011100110010110110110000011100", b"11011110101110101010001101110001"), -- -6.72436e+18 + -1.34614e-21 = -6.72436e+18
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011100110001101101100010000100", b"01111111100000000000000000000000"), -- inf + 1.31585e-21 = inf
	(b"11110100010001100011000101111110", b"00000000000000000000000000000000"),
	(b"11101101000100101010011010011101", b"11110100010001100011001111001001"), -- -6.281e+31 + -2.83664e+27 = -6.28128e+31
	(b"10111011000011100101100101111001", b"00000000000000000000000000000000"),
	(b"11011011100101000110011100011100", b"11011011100101000110011100011100"), -- -0.00217208 + -8.35433e+16 = -8.35433e+16
	(b"01010101100000101100111111001011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.79786e+13 + inf = inf
	(b"00011010011010011000111011000100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.82986e-23 + inf = inf
	(b"00101110001110111111111110000101", b"00000000000000000000000000000000"),
	(b"01101101011101001001000101000001", b"01101101011101001001000101000001"), -- 4.27458e-11 + 4.73062e+27 = 4.73062e+27
	(b"01010100111011010010111101100111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 8.14962e+12 + inf = inf
	(b"00101000010010110000011000101101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.12701e-14 + inf = inf
	(b"00000000000000000000000110001110", b"00000000000000000000000000000000"),
	(b"01000000100101111001101100110110", b"01000000100101111001101100110110"), -- 5.57717e-43 + 4.7377 = 4.7377
	(b"10011111100111100100111101111110", b"00000000000000000000000000000000"),
	(b"10100100010011000010101100111110", b"10100100010011000111101001100110"), -- -6.70471e-20 + -4.42721e-17 = -4.43391e-17
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001011001011110101101001100000", b"10001011001011110101101001100000"), -- -0 + -3.37718e-32 = -3.37718e-32
	(b"10101110100001011011001100010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.07995e-11 + -inf = -inf
	(b"00100011010000111110101111100010", b"00000000000000000000000000000000"),
	(b"00110110101110111010110110000001", b"00110110101110111010110110000001"), -- 1.06209e-17 + 5.59323e-06 = 5.59323e-06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10110001010011001000111111001000", b"00000000000000000000000000000000"),
	(b"11101100010011001000011111011010", b"11101100010011001000011111011010"), -- -2.97676e-09 + -9.8905e+26 = -9.8905e+26
	(b"00101000110110000000011110101100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00101000110110000000011110101100"), -- 2.39841e-14 + 0 = 2.39841e-14
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110101010100000101110001111111", b"11110101010100000101110001111111"), -- -0 + -2.64129e+32 = -2.64129e+32
	(b"00111110010010000000100110010001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0.195349 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01000100101101111110011110000110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1471.24 + inf = inf
	(b"00100000001110000110100101101111", b"00000000000000000000000000000000"),
	(b"01100010011110011001110100101111", b"01100010011110011001110100101111"), -- 1.56203e-19 + 1.15114e+21 = 1.15114e+21
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011011101001010000110111110101", b"00011011101001010000110111110101"), -- 0 + 2.7306e-22 = 2.7306e-22
	(b"01001000101101011011110101000100", b"00000000000000000000000000000000"),
	(b"01011000001010010000100111000001", b"01011000001010010000100111000001"), -- 372202 + 7.43437e+14 = 7.43437e+14
	(b"01010000100010000000000001110011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.82538e+10 + inf = inf
	(b"01000111011101111001101000111101", b"00000000000000000000000000000000"),
	(b"01110000100101111010111110011001", b"01110000100101111010111110011001"), -- 63386.2 + 3.75556e+29 = 3.75556e+29
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110001101001010101011001111101", b"11111111100000000000000000000000"), -- -inf + -1.63743e+30 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100010010000000001101011001011", b"01111111100000000000000000000000"), -- inf + 2.6035e-18 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001100110010100011110011011010", b"01111111100000000000000000000000"), -- inf + 3.11597e-31 = inf
	(b"11001011000110111000100111010000", b"00000000000000000000000000000000"),
	(b"10010011010001111100100111100110", b"11001011000110111000100111010000"), -- -1.01934e+07 + -2.52169e-27 = -1.01934e+07
	(b"10101111101011110101000011111100", b"00000000000000000000000000000000"),
	(b"10111010101000001110010000100010", b"10111010101000001110010000100101"), -- -3.18899e-10 + -0.0012275 = -0.0012275
	(b"10001011010110101000110110111001", b"00000000000000000000000000000000"),
	(b"10101011101111111110101011110100", b"10101011101111111110101011110100"), -- -4.20919e-32 + -1.36366e-12 = -1.36366e-12
	(b"11001001001101111101100001100000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001001001101111101100001100000"), -- -753030 + -0 = -753030
	(b"01101100000011100001101000010011", b"00000000000000000000000000000000"),
	(b"00000001010011101101000111000101", b"01101100000011100001101000010011"), -- 6.87162e+26 + 3.79867e-38 = 6.87162e+26
	(b"01111000100100010011101101100010", b"00000000000000000000000000000000"),
	(b"01001110011001011011010100111011", b"01111000100100010011101101100010"), -- 2.35652e+34 + 9.63465e+08 = 2.35652e+34
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001111100010100110000100111110", b"00001111100010100110000100111110"), -- 0 + 1.36453e-29 = 1.36453e-29
	(b"00011101100010110011000101011011", b"00000000000000000000000000000000"),
	(b"01001011110110110101111100110110", b"01001011110110110101111100110110"), -- 3.6844e-21 + 2.87535e+07 = 2.87535e+07
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100000010101100001100000110101", b"01111111100000000000000000000000"), -- inf + 1.81345e-19 = inf
	(b"10000000000011001100000011101100", b"00000000000000000000000000000000"),
	(b"10011001010101101110111010001111", b"10011001010101101110111010001111"), -- -1.17123e-39 + -1.11117e-23 = -1.11117e-23
	(b"00111000011110110011111011010010", b"00000000000000000000000000000000"),
	(b"00001010100010000011111001100011", b"00111000011110110011111011010010"), -- 5.99016e-05 + 1.31198e-32 = 5.99016e-05
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000100011000001111001010011011", b"01111111100000000000000000000000"), -- inf + 899.791 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11001000110111111110001101111011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -458524 + -inf = -inf
	(b"11000001001000001010010101100101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -10.0404 + -inf = -inf
	(b"01010010100000111000001111101011", b"00000000000000000000000000000000"),
	(b"00000000101001010000100111001110", b"01010010100000111000001111101011"), -- 2.82427e+11 + 1.51564e-38 = 2.82427e+11
	(b"10111001001001110011011010111011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111001001001110011011010111011"), -- -0.000159467 + -0 = -0.000159467
	(b"01000111100110101100101010100100", b"00000000000000000000000000000000"),
	(b"00000001100001100000010100110011", b"01000111100110101100101010100100"), -- 79253.3 + 4.92313e-38 = 79253.3
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001111100011110011100110101101", b"11111111100000000000000000000000"), -- -inf + -4.80584e+09 = -inf
	(b"01001100000001001110011110111011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.48403e+07 + inf = inf
	(b"00101101010101001010110101011100", b"00000000000000000000000000000000"),
	(b"00100011111111011100001001101101", b"00101101010101001010110101111100"), -- 1.20893e-11 + 2.75127e-17 = 1.20893e-11
	(b"01000010111001111001100000111100", b"00000000000000000000000000000000"),
	(b"01111000100100110100010011110111", b"01111000100100110100010011110111"), -- 115.797 + 2.38958e+34 = 2.38958e+34
	(b"11110010110101010110101101101000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110010110101010110101101101000"), -- -8.45442e+30 + -0 = -8.45442e+30
	(b"00111010101000010110110010000001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111010101000010110110010000001"), -- 0.00123157 + 0 = 0.00123157
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000110000101", b"10000000000000000000000110000101"), -- -0 + -5.45105e-43 = -5.45105e-43
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000100010010010001100010101010", b"00000000000000000000000000000000"),
	(b"00111011011011010101011000000001", b"00111011011011010101011000000001"), -- 2.36388e-36 + 0.00362146 = 0.00362146
	(b"01010101000001110111011000100111", b"00000000000000000000000000000000"),
	(b"01100100001011010101110010100110", b"01100100001011010101110010100110"), -- 9.30885e+12 + 1.27919e+22 = 1.27919e+22
	(b"00110101000011100011011010110011", b"00000000000000000000000000000000"),
	(b"00110011110000011100100011000000", b"00110101001001100110111111001011"), -- 5.29787e-07 + 9.02378e-08 = 6.20025e-07
	(b"10000001100110010011000001101110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000001100110010011000001101110"), -- -5.62728e-38 + -0 = -5.62728e-38
	(b"11000001111111111100100010011010", b"00000000000000000000000000000000"),
	(b"11100011100011001111011011101000", b"11100011100011001111011011101000"), -- -31.9729 + -5.20067e+21 = -5.20067e+21
	(b"01001000101011001110101111001101", b"00000000000000000000000000000000"),
	(b"01001010000100000001011010010100", b"01001010001001011011010000001110"), -- 354142 + 2.36074e+06 = 2.71488e+06
	(b"11101011100100110110001110010011", b"00000000000000000000000000000000"),
	(b"10011011100111010010111110010010", b"11101011100100110110001110010011"), -- -3.56365e+26 + -2.60042e-22 = -3.56365e+26
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110101000011100111110011001100", b"00110101000011100111110011001100"), -- 0 + 5.30807e-07 = 5.30807e-07
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001000001100010001101110110001", b"01111111100000000000000000000000"), -- inf + 181359 = inf
	(b"01011000100111111011110111100011", b"00000000000000000000000000000000"),
	(b"01100110001101111111110111001001", b"01100110001101111111110111001001"), -- 1.4051e+15 + 2.17219e+23 = 2.17219e+23
	(b"11111001011010010011111011110100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111001011010010011111011110100"), -- -7.56926e+34 + -0 = -7.56926e+34
	(b"00000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"00000101000110111100000000110111", b"00000101000110111100000000110111"), -- 1.4013e-45 + 7.32337e-36 = 7.32337e-36
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00101001101001010001110100011110", b"00000000000000000000000000000000"),
	(b"00110100000011100011001100000101", b"00110100000011100011001100001010"), -- 7.33252e-14 + 1.32433e-07 = 1.32433e-07
	(b"10100001101011100100101111001100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100001101011100100101111001100"), -- -1.18108e-18 + -0 = -1.18108e-18
	(b"01011000100000001000001001101011", b"00000000000000000000000000000000"),
	(b"00100111111000111110000001110001", b"01011000100000001000001001101011"), -- 1.13038e+15 + 6.32485e-15 = 1.13038e+15
	(b"00101111011100101110010011001110", b"00000000000000000000000000000000"),
	(b"00010001100111110010000101110000", b"00101111011100101110010011001110"), -- 2.20911e-10 + 2.51064e-28 = 2.20911e-10
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00010100110001001101110110110100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.98784e-26 + inf = inf
	(b"10001110000010101010100011010010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10001110000010101010100011010010"), -- -1.70911e-30 + -0 = -1.70911e-30
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000110100100010011001001111010", b"11111111100000000000000000000000"), -- -inf + -18585.2 = -inf
	(b"00010110010011100001101110001110", b"00000000000000000000000000000000"),
	(b"01100110100000111010001111111011", b"01100110100000111010001111111011"), -- 1.66492e-25 + 3.10827e+23 = 3.10827e+23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101001000000101111110111101100", b"00101001000000101111110111101100"), -- 0 + 2.9086e-14 = 2.9086e-14
	(b"00100111001010110011110111110100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.37646e-15 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010000000000000010011001111010", b"01111111100000000000000000000000"), -- inf + 8.60002e+09 = inf
	(b"10111011111000110110111110001000", b"00000000000000000000000000000000"),
	(b"10011001100100111011011010100001", b"10111011111000110110111110001000"), -- -0.00694079 + -1.52732e-23 = -0.00694079
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011100100111001000010010101010", b"10011100100111001000010010101010"), -- -0 + -1.03575e-21 = -1.03575e-21
	(b"11100010001011111110111100111011", b"00000000000000000000000000000000"),
	(b"11010100001111111010100111100111", b"11100010001011111110111100111011"), -- -8.11355e+20 + -3.29276e+12 = -8.11355e+20
	(b"10010001110110011111100110011101", b"00000000000000000000000000000000"),
	(b"11011001101100011111101110011001", b"11011001101100011111101110011001"), -- -3.43904e-28 + -6.26221e+15 = -6.26221e+15
	(b"00011001000010011000000100110101", b"00000000000000000000000000000000"),
	(b"00100011100101101011111010110011", b"00100011100101101011111010110111"), -- 7.10883e-24 + 1.63438e-17 = 1.63438e-17
	(b"00101010000011011111101001110000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.26102e-13 + inf = inf
	(b"10111011000001100000001111100110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0.00204491 + -inf = -inf
	(b"01100110101110100110000001101011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100110101110100110000001101011"), -- 4.40069e+23 + 0 = 4.40069e+23
	(b"11101111001110010110011101111000", b"00000000000000000000000000000000"),
	(b"11110101111111011000010011100100", b"11110101111111011000101010101111"), -- -5.73798e+28 + -6.42747e+32 = -6.42805e+32
	(b"01001010110110100010000011101010", b"00000000000000000000000000000000"),
	(b"01000100100100001101011111000101", b"01001010110110100010100111110111"), -- 7.14764e+06 + 1158.74 = 7.1488e+06
	(b"00011011000111111011101111011110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00011011000111111011101111011110"), -- 1.32129e-22 + 0 = 1.32129e-22
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110110101001111101000101000101", b"01111111100000000000000000000000"), -- inf + 1.70187e+33 = inf
	(b"11000101001010110000100111010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2736.61 + -inf = -inf
	(b"11010011111111100101011110001011", b"00000000000000000000000000000000"),
	(b"10110101111111001111110010011011", b"11010011111111100101011110001011"), -- -2.18478e+12 + -1.8849e-06 = -2.18478e+12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101111101110000011000001001000", b"01101111101110000011000001001000"), -- 0 + 1.14007e+29 = 1.14007e+29
	(b"11001100011010111101101101100000", b"00000000000000000000000000000000"),
	(b"10001000101000111100100110100111", b"11001100011010111101101101100000"), -- -6.18285e+07 + -9.85761e-34 = -6.18285e+07
	(b"10011110011001010111000010011110", b"00000000000000000000000000000000"),
	(b"11000011101101000101111101111100", b"11000011101101000101111101111100"), -- -1.21464e-20 + -360.746 = -360.746
	(b"10100011000011000011100110011101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.60162e-18 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111000001100100010001001011001", b"11111111100000000000000000000000"), -- -inf + -4.24705e-05 = -inf
	(b"00000000000000001100110100101110", b"00000000000000000000000000000000"),
	(b"00011110100010011100000000010111", b"00011110100010011100000000010111"), -- 7.36046e-41 + 1.45849e-20 = 1.45849e-20
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110011110001110001101101101001", b"01111111100000000000000000000000"), -- inf + 9.27165e-08 = inf
	(b"01011001010111001111111010011100", b"00000000000000000000000000000000"),
	(b"00010111010000101000111011000111", b"01011001010111001111111010011100"), -- 3.88778e+15 + 6.2865e-25 = 3.88778e+15
	(b"11011000111101000111111010110110", b"00000000000000000000000000000000"),
	(b"10101010001000101010111100111110", b"11011000111101000111111010110110"), -- -2.1506e+15 + -1.44493e-13 = -2.1506e+15
	(b"01011101110001110010010010001111", b"00000000000000000000000000000000"),
	(b"00110011111111000111010001111111", b"01011101110001110010010010001111"), -- 1.79372e+18 + 1.17559e-07 = 1.79372e+18
	(b"10100010001110100100111110001101", b"00000000000000000000000000000000"),
	(b"11001111001001001011000010010000", b"11001111001001001011000010010000"), -- -2.52498e-18 + -2.76303e+09 = -2.76303e+09
	(b"01011101010011011010110010111011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.26277e+17 + inf = inf
	(b"11001001010011011000001001010000", b"00000000000000000000000000000000"),
	(b"10111110111010001001001111000000", b"11001001010011011000001001010111"), -- -841765 + -0.454252 = -841765
	(b"01100010101000111110101110101011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.5119e+21 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010010000001111100001100010000", b"01111111100000000000000000000000"), -- inf + 1.45773e+11 = inf
	(b"11101000000101110101101000100001", b"00000000000000000000000000000000"),
	(b"11011010100101001010111000100111", b"11101000000101110101101000100001"), -- -2.85896e+24 + -2.09249e+16 = -2.85896e+24
	(b"00100100001001111101001001100010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00100100001001111101001001100010"), -- 3.63906e-17 + 0 = 3.63906e-17
	(b"01100000100101100001011010110011", b"00000000000000000000000000000000"),
	(b"01111111001111000110011111100010", b"01111111001111000110011111100010"), -- 8.65202e+19 + 2.50434e+38 = 2.50434e+38
	(b"10000010000011100011001000000001", b"00000000000000000000000000000000"),
	(b"11011000101100011110100111010100", b"11011000101100011110100111010100"), -- -1.04469e-37 + -1.56494e+15 = -1.56494e+15
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001111000011101111001100111100", b"11001111000011101111001100111100"), -- -0 + -2.39831e+09 = -2.39831e+09
	(b"10101110000011101111110100101101", b"00000000000000000000000000000000"),
	(b"10101111101100110010111001000100", b"10101111110001010000110111101010"), -- -3.25119e-11 + -3.25928e-10 = -3.5844e-10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110100000000010111100110101101", b"11111111100000000000000000000000"), -- -inf + -1.20583e-07 = -inf
	(b"01101110011111111000101101001110", b"00000000000000000000000000000000"),
	(b"00100010110111101010101110000001", b"01101110011111111000101101001110"), -- 1.97718e+28 + 6.03548e-18 = 1.97718e+28
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011101100101000110011011100100", b"01111111100000000000000000000000"), -- inf + 1.33669e+18 = inf
	(b"01001000100011110110001000110001", b"00000000000000000000000000000000"),
	(b"00011001010110101011011111100101", b"01001000100011110110001000110001"), -- 293650 + 1.13075e-23 = 293650
	(b"01101100111000100010101000110110", b"00000000000000000000000000000000"),
	(b"00100100100101110110011111110101", b"01101100111000100010101000110110"), -- 2.18733e+27 + 6.56619e-17 = 2.18733e+27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001111100100011110010001011010", b"10001111100100011110010001011010"), -- -0 + -1.43861e-29 = -1.43861e-29
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11100000010101001110001011010011", b"00000000000000000000000000000000"),
	(b"10000101001010011111011101010001", b"11100000010101001110001011010011"), -- -6.13602e+19 + -7.99177e-36 = -6.13602e+19
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00010000000110011100100101111110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.03292e-29 + inf = inf
	(b"10101010000111110111001101110000", b"00000000000000000000000000000000"),
	(b"11110111000110110001100111110101", b"11110111000110110001100111110101"), -- -1.41621e-13 + -3.14583e+33 = -3.14583e+33
	(b"10001111011111110001100101100101", b"00000000000000000000000000000000"),
	(b"11111101111011100010001110100010", b"11111101111011100010001110100010"), -- -1.25774e-29 + -3.95677e+37 = -3.95677e+37
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110001111011110111001010111000", b"11111111100000000000000000000000"), -- -inf + -6.96886e-09 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101100110110101111101101001101", b"00101100110110101111101101001101"), -- 0 + 6.22383e-12 = 6.22383e-12
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110110001001101100111111010011", b"01111111100000000000000000000000"), -- inf + 8.45836e+32 = inf
	(b"11101000100001100000101101010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.06405e+24 + -inf = -inf
	(b"01000000010001110000111101001111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.11031 + inf = inf
	(b"11111000000011001011111000001100", b"00000000000000000000000000000000"),
	(b"10011100010001100110110110000010", b"11111000000011001011111000001100"), -- -1.14184e+34 + -6.56542e-22 = -1.14184e+34
	(b"00000001100101100010000101000111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.5149e-38 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111000000000000010000100111010", b"11111000000000000010000100111010"), -- -0 + -1.03951e+34 = -1.03951e+34
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001111000000010101010111010000", b"01111111100000000000000000000000"), -- inf + 6.37672e-30 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110110001101011100110101010001", b"01111111100000000000000000000000"), -- inf + 9.21846e+32 = inf
	(b"00101110011000100101011100000110", b"00000000000000000000000000000000"),
	(b"01010110111011011101111111010000", b"01010110111011011101111111010000"), -- 5.14637e-11 + 1.30773e+14 = 1.30773e+14
	(b"01011001010011111000001001100111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.65054e+15 + inf = inf
	(b"01100001000001111011001011111110", b"00000000000000000000000000000000"),
	(b"01101101110111010101100000101011", b"01101101110111010101100000101011"), -- 1.56451e+20 + 8.56285e+27 = 8.56285e+27
	(b"10100001110001011010001100000010", b"00000000000000000000000000000000"),
	(b"11001010101100011001000111001000", b"11001010101100011001000111001000"), -- -1.33924e-18 + -5.8186e+06 = -5.8186e+06
	(b"10101100001111010100100110001101", b"00000000000000000000000000000000"),
	(b"11011110011000010111110001100111", b"11011110011000010111110001100111"), -- -2.68993e-12 + -4.06199e+18 = -4.06199e+18
	(b"01110000001010110110011110101010", b"00000000000000000000000000000000"),
	(b"00110011000001001110111000001110", b"01110000001010110110011110101010"), -- 2.12189e+29 + 3.09502e-08 = 2.12189e+29
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000011010110011", b"00000000000000000000000000000000"),
	(b"01111010001100101101011000110010", b"01111010001100101101011000110010"), -- 2.40323e-42 + 2.32143e+35 = 2.32143e+35
	(b"01110110001011110001001000100101", b"00000000000000000000000000000000"),
	(b"01111011001010111111001100011101", b"01111011001011000001111011100010"), -- 8.87715e+32 + 8.92814e+35 = 8.93701e+35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011001010011000000100000111001", b"11111111100000000000000000000000"), -- -inf + -3.58937e+15 = -inf
	(b"10110100001101111110011110000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.71274e-07 + -inf = -inf
	(b"00111011110001111010010000011000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111011110001111010010000011000"), -- 0.00609256 + 0 = 0.00609256
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01010110110111011111111110001101", b"00000000000000000000000000000000"),
	(b"00110110111100100101111011011000", b"01010110110111011111111110001101"), -- 1.22045e+14 + 7.2232e-06 = 1.22045e+14
	(b"00000000000101111001000000000101", b"00000000000000000000000000000000"),
	(b"01001100001110100111101100111110", b"01001100001110100111101100111110"), -- 2.16388e-39 + 4.8885e+07 = 4.8885e+07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011001100000001110110000101010", b"11111111100000000000000000000000"), -- -inf + -4.53606e+15 = -inf
	(b"01100010101000000101111000000101", b"00000000000000000000000000000000"),
	(b"00110111100010010011110011101001", b"01100010101000000101111000000101"), -- 1.47913e+21 + 1.636e-05 = 1.47913e+21
	(b"01001110010110100111011010100100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001110010110100111011010100100"), -- 9.16302e+08 + 0 = 9.16302e+08
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000101110011", b"11111111100000000000000000000000"), -- -inf + -5.19882e-43 = -inf
	(b"10110100010000000100010110010110", b"00000000000000000000000000000000"),
	(b"10010110111100000010001011011110", b"10110100010000000100010110010110"), -- -1.79067e-07 + -3.87961e-25 = -1.79067e-07
	(b"00000000000000000000000001001010", b"00000000000000000000000000000000"),
	(b"01001111001010101100101000001110", b"01001111001010101100101000001110"), -- 1.03696e-43 + 2.86537e+09 = 2.86537e+09
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111000101000110100111111110111", b"11111000101000110100111111110111"), -- -0 + -2.64989e+34 = -2.64989e+34
	(b"10000000000000000000001101110000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000001110", b"10000000000000000000001101111110"), -- -1.23314e-42 + -1.96182e-44 = -1.25276e-42
	(b"00011000000101010101110101011000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000011011", b"00011000000101010101110101011000"), -- 1.93049e-24 + 3.78351e-44 = 1.93049e-24
	(b"10010000111001110110111110110011", b"00000000000000000000000000000000"),
	(b"10000000000011011000011011010111", b"10010000111001110110111110110011"), -- -9.12855e-29 + -1.24223e-39 = -9.12855e-29
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010101100100101101000110011101", b"01111111100000000000000000000000"), -- inf + 2.01786e+13 = inf
	(b"10111100101011011001101111010000", b"00000000000000000000000000000000"),
	(b"10011001000100100101100100001111", b"10111100101011011001101111010000"), -- -0.0211925 + -7.56601e-24 = -0.0211925
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01010010111011001001111101000101", b"00000000000000000000000000000000"),
	(b"00110111001100011011101001111011", b"01010010111011001001111101000101"), -- 5.08142e+11 + 1.05934e-05 = 5.08142e+11
	(b"10001111010001011111000011010010", b"00000000000000000000000000000000"),
	(b"10100111001101011110000110010111", b"10100111001101011110000110010111"), -- -9.75923e-30 + -2.52411e-15 = -2.52411e-15
	(b"01100000011110111000111110001010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 7.25074e+19 + inf = inf
	(b"00011100001010110111111111000011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000001000", b"00011100001010110111111111000011"), -- 5.67443e-22 + 1.12104e-44 = 5.67443e-22
	(b"10010001110010001100110010000001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10010001110010001100110010000001"), -- -3.16805e-28 + -0 = -3.16805e-28
	(b"11100100100000001001100001000011", b"00000000000000000000000000000000"),
	(b"11100100010000000101111001111011", b"11100100111000001100011110000000"), -- -1.89772e+22 + -1.41943e+22 = -3.31716e+22
	(b"00111110000000111011001001000010", b"00000000000000000000000000000000"),
	(b"01101110110010110010111001111011", b"01101110110010110010111001111011"), -- 0.12861 + 3.14408e+28 = 3.14408e+28
	(b"00110101100011000000001000100110", b"00000000000000000000000000000000"),
	(b"01001101100100011111101111001110", b"01001101100100011111101111001110"), -- 1.04314e-06 + 3.0615e+08 = 3.0615e+08
	(b"11111000000101000111001110101011", b"00000000000000000000000000000000"),
	(b"10100101110010100011101100100001", b"11111000000101000111001110101011"), -- -1.20438e+34 + -3.50815e-16 = -1.20438e+34
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110110010111001100110111101011", b"11110110010111001100110111101011"), -- -0 + -1.11961e+33 = -1.11961e+33
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110010101000111101110010100000", b"11110010101000111101110010100000"), -- -0 + -6.49124e+30 = -6.49124e+30
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001001110010111110011011011110", b"11111111100000000000000000000000"), -- -inf + -4.90876e-33 = -inf
	(b"00101010001011010001101110000001", b"00000000000000000000000000000000"),
	(b"01001101000100011010100110001100", b"01001101000100011010100110001100"), -- 1.5375e-13 + 1.52738e+08 = 1.52738e+08
	(b"01000110111000011110101000000110", b"00000000000000000000000000000000"),
	(b"00010000101010111111000000001101", b"01000110111000011110101000000110"), -- 28917 + 6.78175e-29 = 28917
	(b"01000110010110011001101001011110", b"00000000000000000000000000000000"),
	(b"00111101011011101001010011111110", b"01000110010110011001101010011010"), -- 13926.6 + 0.0582476 = 13926.7
	(b"00101001111101010011101001111000", b"00000000000000000000000000000000"),
	(b"01001001101001001001100111000000", b"01001001101001001001100111000000"), -- 1.08903e-13 + 1.34841e+06 = 1.34841e+06
	(b"11100100110001010000101101111111", b"00000000000000000000000000000000"),
	(b"11001111000001110101010100000111", b"11100100110001010000101101111111"), -- -2.90787e+22 + -2.2705e+09 = -2.90787e+22
	(b"11010001111110010110011011010000", b"00000000000000000000000000000000"),
	(b"10100000100100111111110101011000", b"11010001111110010110011011010000"), -- -1.33896e+11 + -2.50704e-19 = -1.33896e+11
	(b"10010111001100011111011101100101", b"00000000000000000000000000000000"),
	(b"11001100111001111111111010011100", b"11001100111001111111111010011100"), -- -5.7504e-25 + -1.21632e+08 = -1.21632e+08
	(b"00100111111001110110001010001010", b"00000000000000000000000000000000"),
	(b"01010011011110111000011001000011", b"01010011011110111000011001000011"), -- 6.42222e-15 + 1.08029e+12 = 1.08029e+12
	(b"01111101110011110110101000000101", b"00000000000000000000000000000000"),
	(b"01000100110110111110010001101000", b"01111101110011110110101000000101"), -- 3.44626e+37 + 1759.14 = 3.44626e+37
	(b"11010000010110010111110011010111", b"00000000000000000000000000000000"),
	(b"11111110000011111111100001000111", b"11111110000011111111100001000111"), -- -1.45953e+10 + -4.78422e+37 = -4.78422e+37
	(b"10000100000001011110011100100001", b"00000000000000000000000000000000"),
	(b"10010100110100101000101101011100", b"10010100110100101000101101011100"), -- -1.57402e-36 + -2.12595e-26 = -2.12595e-26
	(b"00111110001001011011000100001000", b"00000000000000000000000000000000"),
	(b"01111011000011000011011011000000", b"01111011000011000011011011000000"), -- 0.161808 + 7.28032e+35 = 7.28032e+35
	(b"11100111001000000010000101100110", b"00000000000000000000000000000000"),
	(b"10110001011000000011010110011011", b"11100111001000000010000101100110"), -- -7.56195e+23 + -3.26268e-09 = -7.56195e+23
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010110000100110001011001011101", b"10010110000100110001011001011101"), -- -0 + -1.18816e-25 = -1.18816e-25
	(b"01110101110011010001011100001001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01110101110011010001011100001001"), -- 5.19965e+32 + 0 = 5.19965e+32
	(b"10110011100111001001111000000011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.29306e-08 + -inf = -inf
	(b"00000000000000000000001011100111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000001011100111"), -- 1.04116e-42 + 0 = 1.04116e-42
	(b"11010101101010010110101100111101", b"00000000000000000000000000000000"),
	(b"10011100110110100001001000001100", b"11010101101010010110101100111101"), -- -2.32848e+13 + -1.44307e-21 = -2.32848e+13
	(b"01110000110111001101110000101101", b"00000000000000000000000000000000"),
	(b"00111001101110100101000101110001", b"01110000110111001101110000101101"), -- 5.46823e+29 + 0.000355374 = 5.46823e+29
	(b"01111110110110011111110110000110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.44879e+38 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001111001110111001011000110100", b"11111111100000000000000000000000"), -- -inf + -9.24874e-30 = -inf
	(b"00000011111111100110101001100111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.49532e-36 + inf = inf
	(b"11000010101101101011010000100110", b"00000000000000000000000000000000"),
	(b"10000100101101111111011100100100", b"11000010101101101011010000100110"), -- -91.3519 + -4.32501e-36 = -91.3519
	(b"01001101000111000010100100111101", b"00000000000000000000000000000000"),
	(b"01000001000001100111110101010100", b"01001101000111000010100100111110"), -- 1.63747e+08 + 8.4056 = 1.63747e+08
	(b"10110101011111111010000101010001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -9.52296e-07 + -inf = -inf
	(b"10000011010000000000111000010100", b"00000000000000000000000000000000"),
	(b"11011101010000001100100110001001", b"11011101010000001100100110001001"), -- -5.64399e-37 + -8.68237e+17 = -8.68237e+17
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00010110000001110001110010001001", b"00000000000000000000000000000000"),
	(b"00000110101010111110110011110010", b"00010110000001110001110010001001"), -- 1.09142e-25 + 6.46712e-35 = 1.09142e-25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110110010111111011001000000100", b"11111111100000000000000000000000"), -- -inf + -1.13427e+33 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010011100010011111001010001100", b"01010011100010011111001010001100"), -- 0 + 1.18496e+12 = 1.18496e+12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010111011001110000011010010", b"11111111100000000000000000000000"), -- -inf + -3.33376e+16 = -inf
	(b"11100111100110010000011001011011", b"00000000000000000000000000000000"),
	(b"11010001001110110100001100011110", b"11100111100110010000011001011011"), -- -1.44528e+24 + -5.02678e+10 = -1.44528e+24
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011001011010010010110000001000", b"11111111100000000000000000000000"), -- -inf + -1.20547e-23 = -inf
	(b"00000000000000000010000000100010", b"00000000000000000000000000000000"),
	(b"01101110001010011010110100111111", b"01101110001010011010110100111111"), -- 1.15271e-41 + 1.31281e+28 = 1.31281e+28
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100001111110101101010111001011", b"10100001111110101101010111001011"), -- -0 + -1.69972e-18 = -1.69972e-18
	(b"11001001000110011001010010011000", b"00000000000000000000000000000000"),
	(b"11100111101011110011101100000000", b"11100111101011110011101100000000"), -- -629066 + -1.655e+24 = -1.655e+24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00110100100001110100111101011100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.52035e-07 + inf = inf
	(b"00101101101010110001001010101111", b"00000000000000000000000000000000"),
	(b"01010111010111011101000000111011", b"01010111010111011101000000111011"), -- 1.94487e-11 + 2.43886e+14 = 2.43886e+14
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011110000110011001111110001100", b"11011110000110011001111110001100"), -- -0 + -2.76743e+18 = -2.76743e+18
	(b"00000000000000000000000000000011", b"00000000000000000000000000000000"),
	(b"00110010001011101011010101100101", b"00110010001011101011010101100101"), -- 4.2039e-45 + 1.01694e-08 = 1.01694e-08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00111101110110111010110100011111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111101110110111010110100011111"), -- 0.107264 + 0 = 0.107264
	(b"11000111101110100010011111000000", b"00000000000000000000000000000000"),
	(b"11111000011101101010010100101110", b"11111000011101101010010100101110"), -- -95311.5 + -2.00102e+34 = -2.00102e+34
	(b"00001110011010100001111100010110", b"00000000000000000000000000000000"),
	(b"01011111001001011010110001001010", b"01011111001001011010110001001010"), -- 2.88577e-30 + 1.1938e+19 = 1.1938e+19
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110110100010111111001011010000", b"01110110100010111111001011010000"), -- 0 + 1.41925e+33 = 1.41925e+33
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010111101011100011001111100110", b"11010111101011100011001111100110"), -- -0 + -3.83076e+14 = -3.83076e+14
	(b"01010011010110111101011001010001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.44193e+11 + inf = inf
	(b"01000000010010101110111000110111", b"00000000000000000000000000000000"),
	(b"01001111101101001001011001100100", b"01001111101101001001011001100100"), -- 3.17079 + 6.05951e+09 = 6.05951e+09
	(b"01010001010010011110101101001010", b"00000000000000000000000000000000"),
	(b"01100100100001111101111111111111", b"01100100100001111101111111111111"), -- 5.42022e+10 + 2.00516e+22 = 2.00516e+22
	(b"01101001011100000011100100110010", b"00000000000000000000000000000000"),
	(b"00101001011100101100000110010111", b"01101001011100000011100100110010"), -- 1.81508e+25 + 5.39027e-14 = 1.81508e+25
	(b"00101000001000101010110110100111", b"00000000000000000000000000000000"),
	(b"00111010010010111100111001111110", b"00111010010010111100111001111110"), -- 9.03046e-15 + 0.000777461 = 0.000777461
	(b"00011001000111110011111000011010", b"00000000000000000000000000000000"),
	(b"00100001100101011101110010010101", b"00100001100101011101110011100101"), -- 8.23265e-24 + 1.0155e-18 = 1.01551e-18
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000011100000110010111", b"01000000010000011100000110010111"), -- 0 + 3.02744 = 3.02744
	(b"11000101100101001010000001111000", b"00000000000000000000000000000000"),
	(b"11100001001010010111110101010111", b"11100001001010010111110101010111"), -- -4756.06 + -1.95408e+20 = -1.95408e+20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010000101110011101001110100101", b"10010000101110011101001110100101"), -- -0 + -7.32957e-29 = -7.32957e-29
	(b"11101101110101010101010011011001", b"00000000000000000000000000000000"),
	(b"11100001100001000110100100110110", b"11101101110101010101010011011010"), -- -8.25286e+27 + -3.05319e+20 = -8.25286e+27
	(b"10011111101010100100000010011010", b"00000000000000000000000000000000"),
	(b"10111000100011001010010011111011", b"10111000100011001010010011111011"), -- -7.21047e-20 + -6.70645e-05 = -6.70645e-05
	(b"10011100100111111111010101110011", b"00000000000000000000000000000000"),
	(b"11110110100110100011000100100011", b"11110110100110100011000100100011"), -- -1.05852e-21 + -1.56369e+33 = -1.56369e+33
	(b"11001001010011101111110000101010", b"00000000000000000000000000000000"),
	(b"10001001011000111101001110111001", b"11001001010011101111110000101010"), -- -847811 + -2.74237e-33 = -847811
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100000101100110000010101100001", b"01111111100000000000000000000000"), -- inf + 3.03273e-19 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011101110110111011110010010100", b"11111111100000000000000000000000"), -- -inf + -5.81638e-21 = -inf
	(b"00011011100010010111100000011000", b"00000000000000000000000000000000"),
	(b"01001101000111111011110101001000", b"01001101000111111011110101001000"), -- 2.27424e-22 + 1.67499e+08 = 1.67499e+08
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101101100000011100110110001010", b"01101101100000011100110110001010"), -- 0 + 5.02151e+27 = 5.02151e+27
	(b"11011101000000110010010111011101", b"00000000000000000000000000000000"),
	(b"10111010001110111001000100111000", b"11011101000000110010010111011101"), -- -5.90638e+17 + -0.000715512 = -5.90638e+17
	(b"11000100100101110001101000011111", b"00000000000000000000000000000000"),
	(b"10000101000010011101111011101100", b"11000100100101110001101000011111"), -- -1208.82 + -6.48265e-36 = -1208.82
	(b"11000010110100010111100001000110", b"00000000000000000000000000000000"),
	(b"10011110110000101010001110010000", b"11000010110100010111100001000110"), -- -104.735 + -2.06082e-20 = -104.735
	(b"01100010000010000010001110010101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000011000", b"01100010000010000010001110010101"), -- 6.2783e+20 + 3.36312e-44 = 6.2783e+20
	(b"00001011100000101001110100011100", b"00000000000000000000000000000000"),
	(b"00001011101100100110110101010000", b"00001100000110101000010100110110"), -- 5.03106e-32 + 6.87276e-32 = 1.19038e-31
	(b"11110110010011100101101100110111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110110010011100101101100110111"), -- -1.04635e+33 + -0 = -1.04635e+33
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10100100100010000000000010000011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100100100010000000000010000011"), -- -5.89815e-17 + -0 = -5.89815e-17
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.4013e-45 + -inf = -inf
	(b"10110011101001000110001101110011", b"00000000000000000000000000000000"),
	(b"11100101101111111110100010011111", b"11100101101111111110100010011111"), -- -7.65493e-08 + -1.13283e+23 = -1.13283e+23
	(b"00100101000010000010100010011000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00100101000010000010100010011000"), -- 1.18099e-16 + 0 = 1.18099e-16
	(b"01101101000111100111001101011110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.06488e+27 + inf = inf
	(b"11111001000101001011011101111000", b"00000000000000000000000000000000"),
	(b"11010010100010011111010010001001", b"11111001000101001011011101111000"), -- -4.82613e+34 + -2.96257e+11 = -4.82613e+34
	(b"11100101000101101000101001010001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000101110101", b"11100101000101101000101001010001"), -- -4.44317e+22 + -5.22684e-43 = -4.44317e+22
	(b"00000000001100010010000111011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000001100010010000111011010"), -- 4.51208e-39 + 0 = 4.51208e-39
	(b"00000000010101011011100100000011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000010101011011100100000011"), -- 7.87239e-39 + 0 = 7.87239e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010000000100000111110111011110", b"11111111100000000000000000000000"), -- -inf + -9.69667e+09 = -inf
	(b"00101001111000001101000010100100", b"00000000000000000000000000000000"),
	(b"01010000111000010010001001010011", b"01010000111000010010001001010011"), -- 9.98379e-14 + 3.0217e+10 = 3.0217e+10
	(b"01010101110101000101110001011010", b"00000000000000000000000000000000"),
	(b"01001000101100011011000010111111", b"01010101110101000101110001011010"), -- 2.91866e+13 + 363910 = 2.91866e+13
	(b"00110110100001001101000101000100", b"00000000000000000000000000000000"),
	(b"01110100001011010010110111000111", b"01110100001011010010110111000111"), -- 3.95827e-06 + 5.48826e+31 = 5.48826e+31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000111000101110000100110011011", b"10000111000101110000100110011011"), -- -0 + -1.13628e-34 = -1.13628e-34
	(b"00001011111101000001111111101010", b"00000000000000000000000000000000"),
	(b"01101011111111100000001101100111", b"01101011111111100000001101100111"), -- 9.40334e-32 + 6.14166e+26 = 6.14166e+26
	(b"01010110000111100011001101100100", b"00000000000000000000000000000000"),
	(b"01101100010011001100101111001111", b"01101100010011001100101111001111"), -- 4.34859e+13 + 9.90333e+26 = 9.90333e+26
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11001100110111100100001101010111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001100110111100100001101010111"), -- -1.1653e+08 + -0 = -1.1653e+08
	(b"01101101000101101101011101101110", b"00000000000000000000000000000000"),
	(b"00011010001110010101110010001100", b"01101101000101101101011101101110"), -- 2.9177e+27 + 3.83319e-23 = 2.9177e+27
	(b"00001000011000110100101000011100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.83974e-34 + inf = inf
	(b"11001100110110110110100110101000", b"00000000000000000000000000000000"),
	(b"11111000110001101101110000111001", b"11111000110001101101110000111001"), -- -1.15035e+08 + -3.22669e+34 = -3.22669e+34
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011110010101010100110001101111", b"01011110010101010100110001101111"), -- 0 + 3.84245e+18 = 3.84245e+18
	(b"10010011100101010000000000101000", b"00000000000000000000000000000000"),
	(b"10001101111001100010101110100011", b"10010011100101010000111010001011"), -- -3.7613e-27 + -1.41853e-30 = -3.76272e-27
	(b"01100000101111000001111011011101", b"00000000000000000000000000000000"),
	(b"00011101001111100001001000011100", b"01100000101111000001111011011101"), -- 1.08444e+20 + 2.51557e-21 = 1.08444e+20
	(b"10111111000110100011110111101001", b"00000000000000000000000000000000"),
	(b"11100111101011010000111010111100", b"11100111101011010000111010111100"), -- -0.602507 + -1.63448e+24 = -1.63448e+24
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110001110010011101100111011111", b"11111111100000000000000000000000"), -- -inf + -1.99904e+30 = -inf
	(b"00011100101000101100001111010111", b"00000000000000000000000000000000"),
	(b"01000111101100011000011111111100", b"01000111101100011000011111111100"), -- 1.07709e-21 + 90896 = 90896
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001010000101100110010101111000", b"01001010000101100110010101111000"), -- 0 + 2.46409e+06 = 2.46409e+06
	(b"11100111010101010001000101011101", b"00000000000000000000000000000000"),
	(b"11000011101100100110000001001101", b"11100111010101010001000101011101"), -- -1.00618e+24 + -356.752 = -1.00618e+24
	(b"11110101100100100110000110011000", b"00000000000000000000000000000000"),
	(b"10001100100100000101111100110010", b"11110101100100100110000110011000"), -- -3.7112e+32 + -2.2244e-31 = -3.7112e+32
	(b"11101100000101000011111001011011", b"00000000000000000000000000000000"),
	(b"11100001001000111100001110000111", b"11101100000101000011111001011110"), -- -7.16862e+26 + -1.88807e+20 = -7.16862e+26
	(b"11100101000110001110100010011100", b"00000000000000000000000000000000"),
	(b"11100010111110000000001101101101", b"11100101001000001010100010110111"), -- -4.51307e+22 + -2.28752e+21 = -4.74182e+22
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010001111000101100100000101001", b"00010001111000101100100000101001"), -- 0 + 3.57799e-28 = 3.57799e-28
	(b"11111110000000101100100101001101", b"00000000000000000000000000000000"),
	(b"11000000011111011100101110101110", b"11111110000000101100100101001101"), -- -4.34612e+37 + -3.96556 = -4.34612e+37
	(b"00111001000111110100110111101110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111001000111110100110111101110"), -- 0.000151925 + 0 = 0.000151925
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010100111001010001010001101010", b"01111111100000000000000000000000"), -- inf + 7.87112e+12 = inf
	(b"11010010000110000011001110110110", b"00000000000000000000000000000000"),
	(b"10101101001011010111000101010111", b"11010010000110000011001110110110"), -- -1.63426e+11 + -9.85908e-12 = -1.63426e+11
	(b"10000111110010101011110011110000", b"00000000000000000000000000000000"),
	(b"10110110010000110101111101011100", b"10110110010000110101111101011100"), -- -3.05046e-34 + -2.91128e-06 = -2.91128e-06
	(b"11111101101110100100001110100000", b"00000000000000000000000000000000"),
	(b"10110111110100100011011100101111", b"11111101101110100100001110100000"), -- -3.09484e+37 + -2.50596e-05 = -3.09484e+37
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010010110000010101110110000110", b"01010010110000010101110110000110"), -- 0 + 4.15249e+11 = 4.15249e+11
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000010111001", b"11111111100000000000000000000000"), -- -inf + -2.5924e-43 = -inf
	(b"01011110011010101111100111011001", b"00000000000000000000000000000000"),
	(b"01000101001000010000000100110110", b"01011110011010101111100111011001"), -- 4.23295e+18 + 2576.08 = 4.23295e+18
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111011011000001111110001011010", b"00111011011000001111110001011010"), -- 0 + 0.00343301 = 0.00343301
	(b"11100001101101110010101001111100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.22352e+20 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010110010110010011101001111111", b"01111111100000000000000000000000"), -- inf + 1.75476e-25 = inf
	(b"01100100010111101111110111110111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.64539e+22 + inf = inf
	(b"00100011100010111000111001100011", b"00000000000000000000000000000000"),
	(b"00011100000110101010100011111111", b"00100011100010111000111110011000"), -- 1.51307e-17 + 5.11727e-22 = 1.51312e-17
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10010110000000111011110101011011", b"00000000000000000000000000000000"),
	(b"10001000101101010000011110011010", b"10010110000000111011110101011011"), -- -1.06418e-25 + -1.08953e-33 = -1.06418e-25
	(b"11001101111101110111001011101110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000011010111", b"11001101111101110111001011101110"), -- -5.18938e+08 + -3.01279e-43 = -5.18938e+08
	(b"10010110000110101101100110010101", b"00000000000000000000000000000000"),
	(b"10001010101010000100100100111000", b"10010110000110101101100110010110"), -- -1.25087e-25 + -1.62054e-32 = -1.25087e-25
	(b"01111101001011110001111011101101", b"00000000000000000000000000000000"),
	(b"00000000000001001110001010000111", b"01111101001011110001111011101101"), -- 1.45485e+37 + 4.48605e-40 = 1.45485e+37
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001010101011011001110010101010", b"01111111100000000000000000000000"), -- inf + 5.68892e+06 = inf
	(b"00000101111111101010110010100110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000101111111101010110010100110"), -- 2.39495e-35 + 0 = 2.39495e-35
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001001100111100000100101001000", b"00001001100111100000100101001000"), -- 0 + 3.80458e-33 = 3.80458e-33
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011011101011110111010010001000", b"01111111100000000000000000000000"), -- inf + 9.87725e+16 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010100101100011000000001111010", b"11111111100000000000000000000000"), -- -inf + -1.79231e-26 = -inf
	(b"11001101110000011101001100010001", b"00000000000000000000000000000000"),
	(b"11010101010000100100110001010110", b"11010101010000100100110111011010"), -- -4.06479e+08 + -1.33521e+13 = -1.33525e+13
	(b"00001111001011110010101101001111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 8.63651e-30 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010001001110001101100000011010", b"11010001001110001101100000011010"), -- -0 + -4.96187e+10 = -4.96187e+10
	(b"01010110011001100110110001010111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.33382e+13 + inf = inf
	(b"11000000001111100100111000010011", b"00000000000000000000000000000000"),
	(b"11011101000001000001010001001000", b"11011101000001000001010001001000"), -- -2.97352 + -5.94832e+17 = -5.94832e+17
	(b"11110101111000101100000010100111", b"00000000000000000000000000000000"),
	(b"11101000001010000001111101010100", b"11110101111000101100000010100111"), -- -5.74886e+32 + -3.17574e+24 = -5.74886e+32
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101100100010111100011000110111", b"01101100100010111100011000110111"), -- 0 + 1.35181e+27 = 1.35181e+27
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010100000110101000000111100101", b"00010100000110101000000111100101"), -- 0 + 7.80063e-27 = 7.80063e-27
	(b"11011100111111010101110111110111", b"00000000000000000000000000000000"),
	(b"10010110101001110010010011011110", b"11011100111111010101110111110111"), -- -5.70532e+17 + -2.70036e-25 = -5.70532e+17
	(b"00111000100011111101000111010001", b"00000000000000000000000000000000"),
	(b"00001000110111100010110100110000", b"00111000100011111101000111010001"), -- 6.85785e-05 + 1.33718e-33 = 6.85785e-05
	(b"11001001000010101111010011100000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -569166 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110010100011111011001100101101", b"10110010100011111011001100101101"), -- -0 + -1.67289e-08 = -1.67289e-08
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000001", b"00000000000000000000000000000001"), -- 0 + 1.4013e-45 = 1.4013e-45
	(b"11010111111100001001001111011000", b"00000000000000000000000000000000"),
	(b"10000000100010110000011001100100", b"11010111111100001001001111011000"), -- -5.29036e+14 + -1.27674e-38 = -5.29036e+14
	(b"11000111101111110100101001000111", b"00000000000000000000000000000000"),
	(b"10010010000100010101101000000000", b"11000111101111110100101001000111"), -- -97940.6 + -4.58649e-28 = -97940.6
	(b"10010011100001001111000111110110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10010011100001001111000111110110"), -- -3.35601e-27 + -0 = -3.35601e-27
	(b"11101110100111010010111110110011", b"00000000000000000000000000000000"),
	(b"10101000000100000010011000001111", b"11101110100111010010111110110011"), -- -2.43234e+28 + -8.00186e-15 = -2.43234e+28
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10001010001010100110100000001011", b"00000000000000000000000000000000"),
	(b"11010001110011010010010000100110", b"11010001110011010010010000100110"), -- -8.20477e-33 + -1.10134e+11 = -1.10134e+11
	(b"00100100010110001000100001111100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.69531e-17 + inf = inf
	(b"11000011000010010100010111000111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -137.273 + -inf = -inf
	(b"10110000010100111111101111010000", b"00000000000000000000000000000000"),
	(b"10110111011110000110001111111001", b"10110111011110000110011101001001"), -- -7.71192e-10 + -1.48052e-05 = -1.4806e-05
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01010111100011011000110010110111", b"00000000000000000000000000000000"),
	(b"00011000001110010111101010110010", b"01010111100011011000110010110111"), -- 3.11271e+14 + 2.39726e-24 = 3.11271e+14
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011111100110110011000011", b"11000000011111100110110011000011"), -- -0 + -3.97539 = -3.97539
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11010010101010101011111101011101", b"00000000000000000000000000000000"),
	(b"10101011110111001011011100100001", b"11010010101010101011111101011101"), -- -3.66677e+11 + -1.56828e-12 = -3.66677e+11
	(b"10100000101101101000011111110000", b"00000000000000000000000000000000"),
	(b"10010101100000000000101101001111", b"10100000101101101000011111110010"), -- -3.0922e-19 + -5.17166e-26 = -3.0922e-19
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010111101101110100010111000010", b"10010111101101110100010111000010"), -- -0 + -1.18437e-24 = -1.18437e-24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"01100001100100001001010010010011", b"01100001100100001001010010010011"), -- 1.4013e-45 + 3.3338e+20 = 3.3338e+20
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010011101011101010101101111001", b"00010011101011101010101101111001"), -- 0 + 4.40929e-27 = 4.40929e-27
	(b"01011111010000110001111101100110", b"00000000000000000000000000000000"),
	(b"00010011111111001101100010101001", b"01011111010000110001111101100110"), -- 1.40601e+19 + 6.38274e-27 = 1.40601e+19
	(b"01010010111010100111001101110001", b"00000000000000000000000000000000"),
	(b"00010101010011000101000110010110", b"01010010111010100111001101110001"), -- 5.0348e+11 + 4.12618e-26 = 5.0348e+11
	(b"00010011000001100011010011011100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.69392e-27 + inf = inf
	(b"00000000000000001001010111111001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.38001e-41 + inf = inf
	(b"00111000010101000011001101101101", b"00000000000000000000000000000000"),
	(b"00000101100101100111100000000110", b"00111000010101000011001101101101"), -- 5.05926e-05 + 1.415e-35 = 5.05926e-05
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010011101000011001100110", b"01000010010011101000011001100110"), -- 0 + 51.6312 = 51.6312
	(b"00101101000100111110011001010010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 8.40712e-12 + inf = inf
	(b"10001000000000101110100101001100", b"00000000000000000000000000000000"),
	(b"10110000101001111000001010111111", b"10110000101001111000001010111111"), -- -3.93947e-34 + -1.2188e-09 = -1.2188e-09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100000111110100101001", b"01111111100000000000000000000000"), -- inf + 2.75764 = inf
	(b"11001100111100010100100101101100", b"00000000000000000000000000000000"),
	(b"10111000001000000000110110010100", b"11001100111100010100100101101100"), -- -1.26504e+08 + -3.81596e-05 = -1.26504e+08
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011110111000000010000000011111", b"01111111100000000000000000000000"), -- inf + 2.37302e-20 = inf
	(b"01111110111000110010111111000001", b"00000000000000000000000000000000"),
	(b"00100111000001101100010010101101", b"01111110111000110010111111000001"), -- 1.50991e+38 + 1.87029e-15 = 1.50991e+38
	(b"10110011010000010000000101111010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110011010000010000000101111010"), -- -4.49377e-08 + -0 = -4.49377e-08
	(b"00000000000000000000111010110111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.27869e-42 + inf = inf
	(b"01110000101011000111100101001011", b"00000000000000000000000000000000"),
	(b"01111010100110110011011101000010", b"01111010100110110011011101001101"), -- 4.27024e+29 + 4.02963e+35 = 4.02964e+35
	(b"11010100000001010101000111001110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.29041e+12 + -inf = -inf
	(b"11011001101110001011100100010110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.49936e+15 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011001000010100010101111100110", b"01011001000010100010101111100110"), -- 0 + 2.43074e+15 = 2.43074e+15
	(b"10101011010011000011100111000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.25555e-13 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100001101100011100110101100001", b"00100001101100011100110101100001"), -- 0 + 1.20483e-18 = 1.20483e-18
	(b"11110011101000101111010001111011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.58213e+31 + -inf = -inf
	(b"01111110101011100110101000101010", b"00000000000000000000000000000000"),
	(b"00111000000101100100101000011111", b"01111110101011100110101000101010"), -- 1.15918e+38 + 3.58318e-05 = 1.15918e+38
	(b"01011011000001001101110011011101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01011011000001001101110011011101"), -- 3.73975e+16 + 0 = 3.73975e+16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001000111101110011001001011110", b"11111111100000000000000000000000"), -- -inf + -1.48776e-33 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001011101010001100110100011001", b"01111111100000000000000000000000"), -- inf + 6.50198e-32 = inf
	(b"11100011110001100111110010110110", b"00000000000000000000000000000000"),
	(b"10000000000000000000100010100010", b"11100011110001100111110010110110"), -- -7.32288e+21 + -3.09687e-42 = -7.32288e+21
	(b"10111000001000010011100011000101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.84383e-05 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100010101000101000011010011100", b"10100010101000101000011010011100"), -- -0 + -4.40527e-18 = -4.40527e-18
	(b"10011011101011010101110101100000", b"00000000000000000000000000000000"),
	(b"11001100101110111011011010100000", b"11001100101110111011011010100000"), -- -2.86808e-22 + -9.84159e+07 = -9.84159e+07
	(b"00010011100001010111110001000000", b"00000000000000000000000000000000"),
	(b"01001110101010001001111100101111", b"01001110101010001001111100101111"), -- 3.36964e-27 + 1.4145e+09 = 1.4145e+09
	(b"00111110001101000001110011010111", b"00000000000000000000000000000000"),
	(b"01001011100100100101101101011111", b"01001011100100100101101101011111"), -- 0.175891 + 1.91833e+07 = 1.91833e+07
	(b"11111100000000100110111110110010", b"00000000000000000000000000000000"),
	(b"10111101110011010100111100101001", b"11111100000000100110111110110010"), -- -2.70906e+36 + -0.100249 = -2.70906e+36
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011000001110110100001110000101", b"11111111100000000000000000000000"), -- -inf + -2.42033e-24 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01000000110100010001100010110100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.53427 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110000110000000000001100", b"10111110110000110000000000001100"), -- -0 + -0.38086 = -0.38086
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000100111110000111111", b"00000000000000100111110000111111"), -- 0 + 2.28242e-40 = 2.28242e-40
	(b"11010111000000000010100001110011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.40911e+14 + -inf = -inf
	(b"10110110101101111010011101010001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.4733e-06 + -inf = -inf
	(b"11011101001001010010101100100010", b"00000000000000000000000000000000"),
	(b"11110100010110101010010101111111", b"11110100010110101010010101111111"), -- -7.43853e+17 + -6.92918e+31 = -6.92918e+31
	(b"01001111010100111000001111010101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001111010100111000001111010101"), -- 3.54863e+09 + 0 = 3.54863e+09
	(b"00110110011011000101001100000111", b"00000000000000000000000000000000"),
	(b"00011101100101111100011000100101", b"00110110011011000101001100000111"), -- 3.52151e-06 + 4.01742e-21 = 3.52151e-06
	(b"01010101100101010111001100010011", b"00000000000000000000000000000000"),
	(b"01000001100100101010100000011010", b"01010101100101010111001100010011"), -- 2.05402e+13 + 18.3321 = 2.05402e+13
	(b"00100101111011010010000110001110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.11357e-16 + inf = inf
	(b"10000010001111111100111100111101", b"00000000000000000000000000000000"),
	(b"10100001110111110100110001011111", b"10100001110111110100110001011111"), -- -1.40919e-37 + -1.51313e-18 = -1.51313e-18
	(b"10000011110011110001000001110001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.21701e-36 + -inf = -inf
	(b"00000000000000001001010000101010", b"00000000000000000000000000000000"),
	(b"00010111110100101101010100101101", b"00010111110100101101010100101101"), -- 5.31513e-41 + 1.36247e-24 = 1.36247e-24
	(b"11100010100011011101011111110101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.30828e+21 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010010101111100010000011000000", b"00010010101111100010000011000000"), -- 0 + 1.19988e-27 = 1.19988e-27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000010100000101010101", b"10000000000000010100000101010101"), -- -0 + -1.15272e-40 = -1.15272e-40
	(b"00100111101001111011111100011100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00100111101001111011111100011100"), -- 4.6559e-15 + 0 = 4.6559e-15
	(b"01100111100101000110000010010111", b"00000000000000000000000000000000"),
	(b"00111101011011100110000100001111", b"01100111100101000110000010010111"), -- 1.40138e+24 + 0.058198 = 1.40138e+24
	(b"00111001100010101010100110101000", b"00000000000000000000000000000000"),
	(b"00010001110001011001100011000110", b"00111001100010101010100110101000"), -- 0.000264478 + 3.11753e-28 = 0.000264478
	(b"11110000010001000111010000101010", b"00000000000000000000000000000000"),
	(b"10010101100011000100110011110001", b"11110000010001000111010000101010"), -- -2.43198e+29 + -5.66669e-26 = -2.43198e+29
	(b"00111001110001101111010100011111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0.000379481 + inf = inf
	(b"10100100100110011010100011011100", b"00000000000000000000000000000000"),
	(b"10011110110001110110100100011001", b"10100100100110011011010101010011"), -- -6.66392e-17 + -2.11134e-20 = -6.66603e-17
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111001100100001100111001111000", b"01111111100000000000000000000000"), -- inf + 0.000276197 = inf
	(b"10110110010010100111011010010110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000101001111", b"10110110010010100111011010010110"), -- -3.01694e-06 + -4.69435e-43 = -3.01694e-06
	(b"10101111010111011001100001111000", b"00000000000000000000000000000000"),
	(b"10001101100100011001011001001001", b"10101111010111011001100001111000"), -- -2.0154e-10 + -8.97249e-31 = -2.0154e-10
	(b"00101111101100011000110101000101", b"00000000000000000000000000000000"),
	(b"00100100100011111010010100000001", b"00101111101100011000110101000111"), -- 3.22965e-10 + 6.22959e-17 = 3.22965e-10
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11010110010101111101100011010111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.93316e+13 + -inf = -inf
	(b"10000000000000000000000001010001", b"00000000000000000000000000000000"),
	(b"10000010010101100110000010110001", b"10000010010101100110000010111011"), -- -1.13505e-43 + -1.575e-37 = -1.575e-37
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111011000101000001001110011000", b"11111111100000000000000000000000"), -- -inf + -0.00225947 = -inf
	(b"01101111001110000110000011110000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.70624e+28 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000101000000011111111001100111", b"11111111100000000000000000000000"), -- -inf + -2079.9 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011110110110000110110001011", b"11111111100000000000000000000000"), -- -inf + -2.87117e+07 = -inf
	(b"11010001000011100001000001110110", b"00000000000000000000000000000000"),
	(b"10000000000011001101101001101110", b"11010001000011100001000001110110"), -- -3.81351e+10 + -1.18038e-39 = -3.81351e+10
	(b"10011001010001111110010011101101", b"00000000000000000000000000000000"),
	(b"10111001101010100111011101001101", b"10111001101010100111011101001101"), -- -1.03343e-23 + -0.000325138 = -0.000325138
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110001010110001101001110101000", b"01111111100000000000000000000000"), -- inf + 3.15524e-09 = inf
	(b"10010101110110100110111100000111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.82247e-26 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010000110010010100010011", b"11111111100000000000000000000000"), -- -inf + -0.190571 = -inf
	(b"11101001011000101010111011001100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11101001011000101010111011001100"), -- -1.71277e+25 + -0 = -1.71277e+25
	(b"11001000101010010000110110011101", b"00000000000000000000000000000000"),
	(b"10100010101011001101110000000010", b"11001000101010010000110110011101"), -- -346221 + -4.68536e-18 = -346221
	(b"01011111011101010010001101111000", b"00000000000000000000000000000000"),
	(b"01000001011000001110001000101000", b"01011111011101010010001101111000"), -- 1.76641e+19 + 14.0552 = 1.76641e+19
	(b"01010001101100101001011110011001", b"00000000000000000000000000000000"),
	(b"01100001100010101001110100011010", b"01100001100010101001110100011010"), -- 9.58809e+10 + 3.19621e+20 = 3.19621e+20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010000110011010000111010010001", b"11010000110011010000111010010001"), -- -0 + -2.75223e+10 = -2.75223e+10
	(b"01110101011010110010101001110111", b"00000000000000000000000000000000"),
	(b"00101011000010011001001110111111", b"01110101011010110010101001110111"), -- 2.98108e+32 + 4.88772e-13 = 2.98108e+32
	(b"00000100110111101000111100100000", b"00000000000000000000000000000000"),
	(b"01101101000000011011010101100010", b"01101101000000011011010101100010"), -- 5.23234e-36 + 2.50893e+27 = 2.50893e+27
	(b"10011000010001011111010010111100", b"00000000000000000000000000000000"),
	(b"10110011110100010010000000000000", b"10110011110100010010000000000000"), -- -2.55852e-24 + -9.73814e-08 = -9.73814e-08
	(b"10010111000100010110111111100111", b"00000000000000000000000000000000"),
	(b"10100011110010011110010000110101", b"10100011110010011110010000110101"), -- -4.69933e-25 + -2.18891e-17 = -2.18891e-17
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100110011010100100011000110111", b"01111111100000000000000000000000"), -- inf + 2.76582e+23 = inf
	(b"00000000010100111011010101001100", b"00000000000000000000000000000000"),
	(b"00111010100100101101010011111011", b"00111010100100101101010011111011"), -- 7.68738e-39 + 0.00112024 = 0.00112024
	(b"00011001001101101101100110010100", b"00000000000000000000000000000000"),
	(b"00100101100001100000010101111000", b"00100101100001100000010101111000"), -- 9.45312e-24 + 2.3249e-16 = 2.3249e-16
	(b"11000100010011100010111011010001", b"00000000000000000000000000000000"),
	(b"10010011010101001001110100101000", b"11000100010011100010111011010001"), -- -824.732 + -2.68356e-27 = -824.732
	(b"11101111111101001101001011000010", b"00000000000000000000000000000000"),
	(b"10011100000110100111010100111001", b"11101111111101001101001011000010"), -- -1.51538e+29 + -5.11058e-22 = -1.51538e+29
	(b"11110001101000011011111010011011", b"00000000000000000000000000000000"),
	(b"11101111111101011110100010110110", b"11110001101100010001110100100110"), -- -1.60184e+30 + -1.5221e+29 = -1.75405e+30
	(b"00110000110101000100110110101100", b"00000000000000000000000000000000"),
	(b"00110110001011101111011101111000", b"00110110001011110001001000000010"), -- 1.54471e-09 + 2.60721e-06 = 2.60875e-06
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000010101100011", b"00000000000000000000000000000000"),
	(b"01111000111000110111001011101000", b"01111000111000110111001011101000"), -- 1.93239e-42 + 3.69057e+34 = 3.69057e+34
	(b"00011101111100010011111111101101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.38583e-21 + inf = inf
	(b"11101111110111111110101111101000", b"00000000000000000000000000000000"),
	(b"10110111100001101010000000000111", b"11101111110111111110101111101000"), -- -1.38601e+29 + -1.60486e-05 = -1.38601e+29
	(b"11000001011000011100111110111000", b"00000000000000000000000000000000"),
	(b"10000001001011010111111100001110", b"11000001011000011100111110111000"), -- -14.1132 + -3.18662e-38 = -14.1132
	(b"00011000011100001011010101011000", b"00000000000000000000000000000000"),
	(b"00100111110101111011111000100101", b"00100111110101111011111000100101"), -- 3.11108e-24 + 5.98806e-15 = 5.98806e-15
	(b"00011011001010001010101111100001", b"00000000000000000000000000000000"),
	(b"00011011011110111100111101011110", b"00011011110100100011110110100000"), -- 1.39522e-22 + 2.08292e-22 = 3.47814e-22
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01010010101000100111010011101101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.48873e+11 + inf = inf
	(b"01011000100001011010011110111011", b"00000000000000000000000000000000"),
	(b"01001101101000010110101100001100", b"01011000100001011010011110111110"), -- 1.17564e+15 + 3.38518e+08 = 1.17564e+15
	(b"00110011101001011011001111010011", b"00000000000000000000000000000000"),
	(b"01100100101110100011100111110000", b"01100100101110100011100111110000"), -- 7.71612e-08 + 2.74822e+22 = 2.74822e+22
	(b"00001101100000010011101111110010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00001101100000010011101111110010"), -- 7.96467e-31 + 0 = 7.96467e-31
	(b"00011010000010010111111001101100", b"00000000000000000000000000000000"),
	(b"01111110010110110011111001000101", b"01111110010110110011111001000101"), -- 2.84331e-23 + 7.28561e+37 = 7.28561e+37
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000011101001111000011111100111", b"01111111100000000000000000000000"), -- inf + 335.062 = inf
	(b"11100100101010100011010010000101", b"00000000000000000000000000000000"),
	(b"11101011011000010101110000011001", b"11101011011000010110000101101011"), -- -2.51178e+22 + -2.72443e+26 = -2.72468e+26
	(b"00111000010000111010000101111000", b"00000000000000000000000000000000"),
	(b"01011100100100010011101000111111", b"01011100100100010011101000111111"), -- 4.6642e-05 + 3.27023e+17 = 3.27023e+17
	(b"10100000110000110101101111111111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.30952e-19 + -inf = -inf
	(b"11110101001011001010100101000011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.18874e+32 + -inf = -inf
	(b"01001111101011101101101100011001", b"00000000000000000000000000000000"),
	(b"00010111010111101010010000111110", b"01001111101011101101101100011001"), -- 5.86719e+09 + 7.19394e-25 = 5.86719e+09
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010010101001010001111010101111", b"10010010101001010001111010101111"), -- -0 + -1.04205e-27 = -1.04205e-27
	(b"01000000001000110101010000101110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000000001000110101010000101110"), -- 2.55201 + 0 = 2.55201
	(b"00000000000000000000000000101001", b"00000000000000000000000000000000"),
	(b"00011001111111100101010100101011", b"00011001111111100101010100101011"), -- 5.74532e-44 + 2.62974e-23 = 2.62974e-23
	(b"00011011000110110111000011111010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00011011000110110111000011111010"), -- 1.28578e-22 + 0 = 1.28578e-22
	(b"01010100000100011111001010100001", b"00000000000000000000000000000000"),
	(b"01000100001101010010100110101000", b"01010100000100011111001010100001"), -- 2.50736e+12 + 724.651 = 2.50736e+12
	(b"00011101000000110011011001000001", b"00000000000000000000000000000000"),
	(b"00001100101101011010111110101110", b"00011101000000110011011001000001"), -- 1.73658e-21 + 2.79932e-31 = 1.73658e-21
	(b"10011110000111110000010111100010", b"00000000000000000000000000000000"),
	(b"11110110000010000000110111101100", b"11110110000010000000110111101100"), -- -8.41861e-21 + -6.89878e+32 = -6.89878e+32
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100011111011101111101001001010", b"01111111100000000000000000000000"), -- inf + 2.591e-17 = inf
	(b"10110111000001101111101010010101", b"00000000000000000000000000000000"),
	(b"11010100110111001101001100000001", b"11010100110111001101001100000001"), -- -8.04537e-06 + -7.58746e+12 = -7.58746e+12
	(b"10011011000010001100011101100010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.13141e-22 + -inf = -inf
	(b"11100111001100100011100011001101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.41629e+23 + -inf = -inf
	(b"00000000000000000000000001101001", b"00000000000000000000000000000000"),
	(b"00100000110111101111110001011000", b"00100000110111101111110001011000"), -- 1.47136e-43 + 3.77752e-19 = 3.77752e-19
	(b"10101110000001111000001001001001", b"00000000000000000000000000000000"),
	(b"11111100010000101011110010101000", b"11111100010000101011110010101000"), -- -3.08112e-11 + -4.04453e+36 = -4.04453e+36
	(b"00010110011110101101001000000110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00010110011110101101001000000110"), -- 2.02611e-25 + 0 = 2.02611e-25
	(b"00011100100011100010110010011101", b"00000000000000000000000000000000"),
	(b"01100110101000010101110111101110", b"01100110101000010101110111101110"), -- 9.4083e-22 + 3.81017e+23 = 3.81017e+23
	(b"01000010011001101101000011111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000010011001101101000011111011"), -- 57.7041 + 0 = 57.7041
	(b"00000001110100101011100111100110", b"00000000000000000000000000000000"),
	(b"01100010111010111100011100000111", b"01100010111010111100011100000111"), -- 7.74086e-38 + 2.17466e+21 = 2.17466e+21
	(b"01110011001010110000000010100010", b"00000000000000000000000000000000"),
	(b"01001010010101111000001011110101", b"01110011001010110000000010100010"), -- 1.35482e+31 + 3.53094e+06 = 1.35482e+31
	(b"01010100001000001011111010101001", b"00000000000000000000000000000000"),
	(b"01001011100100000000101010111111", b"01010100001000001011111011110001"), -- 2.76157e+12 + 1.88799e+07 = 2.76159e+12
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000110", b"00000000000000000000000000000110"), -- 0 + 8.40779e-45 = 8.40779e-45
	(b"10111100011111111111101110110000", b"00000000000000000000000000000000"),
	(b"10011101100110000010011100110011", b"10111100011111111111101110110000"), -- -0.015624 + -4.02746e-21 = -0.015624
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011101111110001011110111100000", b"01111111100000000000000000000000"), -- inf + 6.58414e-21 = inf
	(b"00011111010011101110011101001010", b"00000000000000000000000000000000"),
	(b"01011101010101101001010101110001", b"01011101010101101001010101110001"), -- 4.38135e-20 + 9.66399e+17 = 9.66399e+17
	(b"01010001010011101100000100100000", b"00000000000000000000000000000000"),
	(b"00010011011001011010110011111001", b"01010001010011101100000100100000"), -- 5.55002e+10 + 2.89891e-27 = 5.55002e+10
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01011100010110111100001111101010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.47434e+17 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110100100010101100001111001111", b"01111111100000000000000000000000"), -- inf + 8.79527e+31 = inf
	(b"11101100001101011100110100001100", b"00000000000000000000000000000000"),
	(b"10000111010110100101001101111101", b"11101100001101011100110100001100"), -- -8.79136e+26 + -1.6425e-34 = -8.79136e+26
	(b"11101101010000101101000000011010", b"00000000000000000000000000000000"),
	(b"11110001100010000011101010000010", b"11110001100010001001101111101010"), -- -3.76823e+27 + -1.34914e+30 = -1.35291e+30
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000001"), -- -1.4013e-45 + -0 = -1.4013e-45

	(b"11101111111101010111111100100011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11101111111101010111111100100011"), -- -1.51955e+29 + -0 = -1.51955e+29
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01000010100011110010011110011010", b"00000000000000000000000000000000"),
	(b"01100100011010001111100010001101", b"01100100011010001111100010001101"), -- 71.5773 + 1.71902e+22 = 1.71902e+22
	(b"00000011000001110011011101011100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.97365e-37 + inf = inf
	(b"10100001001100011011010110101001", b"00000000000000000000000000000000"),
	(b"10000011000110111011111100111010", b"10100001001100011011010110101001"), -- -6.02104e-19 + -4.57699e-37 = -6.02104e-19
	(b"00110010101101010100101111010000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.11056e-08 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011001010101100100010100111101", b"11011001010101100100010100111101"), -- -0 + -3.76949e+15 = -3.76949e+15
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110011101101000001101111111110", b"11111111100000000000000000000000"), -- -inf + -2.85395e+31 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001000110111000001011100", b"00111111001000110111000001011100"), -- 0 + 0.638433 = 0.638433
	(b"00011100110011010000000101011000", b"00000000000000000000000000000000"),
	(b"01010110010011110101111111101001", b"01010110010011110101111111101001"), -- 1.35661e-21 + 5.70027e+13 = 5.70027e+13
	(b"11011010101000111110010101101101", b"00000000000000000000000000000000"),
	(b"10011011110101111110110000010111", b"11011010101000111110010101101101"), -- -2.30663e+16 + -3.57213e-22 = -2.30663e+16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101001100011111110001000001010", b"11111111100000000000000000000000"), -- -inf + -6.38969e-14 = -inf
	(b"10000000000000000000010111111001", b"00000000000000000000000000000000"),
	(b"11111010100101000011110000001111", b"11111010100101000011110000001111"), -- -2.14259e-42 + -3.84839e+35 = -3.84839e+35
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101110001100101110101011111011", b"11101110001100101110101011111011"), -- -0 + -1.38431e+28 = -1.38431e+28
	(b"01101011001100010110101010101110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.14484e+26 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00110101110101000101111111011111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.58231e-06 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100001010000110010011001011011", b"11100001010000110010011001011011"), -- -0 + -2.24992e+20 = -2.24992e+20
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000101010000100101101001110101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -9.13845e-36 + -inf = -inf
	(b"00000000000000001011101101001100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.71895e-41 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000100110001", b"11111111100000000000000000000000"), -- -inf + -4.27396e-43 = -inf
	(b"10010000101001001101100000110010", b"00000000000000000000000000000000"),
	(b"11011100000110110100110001110110", b"11011100000110110100110001110110"), -- -6.50197e-29 + -1.74851e+17 = -1.74851e+17
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01000101001111101001110111011011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000101001111101001110111011011"), -- 3049.87 + 0 = 3049.87
	(b"10101001011011000101000000110011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.24721e-14 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011101101101010101000111110110", b"10011101101101010101000111110110"), -- -0 + -4.7995e-21 = -4.7995e-21
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000001010000011000111100", b"00000000000001010000011000111100"), -- 0 + 4.61414e-40 = 4.61414e-40
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111010011010111010100110110011", b"01111111100000000000000000000000"), -- inf + 0.000898983 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10001010000000100000010011001011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.26017e-33 + -inf = -inf
	(b"01101111000101001000111011000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101111000101001000111011000000"), -- 4.59764e+28 + 0 = 4.59764e+28
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101011110011010000111011101101", b"11101011110011010000111011101101"), -- -0 + -4.95801e+26 = -4.95801e+26
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011000100010100101000010101001", b"01111111100000000000000000000000"), -- inf + 3.57536e-24 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010011001011100000011011100100", b"00010011001011100000011011100100"), -- 0 + 2.19653e-27 = 2.19653e-27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11110110001111100000011111000111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110110001111100000011111000111"), -- -9.63569e+32 + -0 = -9.63569e+32
	(b"00101011110111101111110100101001", b"00000000000000000000000000000000"),
	(b"00100101101111011111100111101011", b"00101011110111110000100100001001"), -- 1.58443e-12 + 3.29556e-16 = 1.58476e-12
	(b"10110101101111111001011100010000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110101101111111001011100010000"), -- -1.42746e-06 + -0 = -1.42746e-06
	(b"10111010101100110010110011001110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111010101100110010110011001110"), -- -0.001367 + -0 = -0.001367
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01110101010010111011110000101100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.58265e+32 + inf = inf
	(b"00011011101010110001100001110010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.83054e-22 + inf = inf
	(b"10011001100000001001000110100001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10011001100000001001000110100001"), -- -1.32937e-23 + -0 = -1.32937e-23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000100111001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.38606e-43 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11100011000011001001011101000110", b"00000000000000000000000000000000"),
	(b"11101001000011001010101110101011", b"11101001000011001011010001110100"), -- -2.59344e+21 + -1.06288e+25 = -1.06314e+25
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10111111011010011011111111010110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111011010011011111111010110"), -- -0.913083 + -0 = -0.913083
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001111100101001101000001111", b"11111111100000000000000000000000"), -- -inf + -3.66609e+25 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11001101001100000101000101100110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.84883e+08 + -inf = -inf
	(b"11110111101100010101001111000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110111101100010101001111000000"), -- -7.19324e+33 + -0 = -7.19324e+33
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000100010001010100001111111010", b"01000100010001010100001111111010"), -- 0 + 789.062 = 789.062
	(b"00000000000000000000011000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000011000000000"), -- 2.15239e-42 + 0 = 2.15239e-42
	(b"01110101110101100111000000010100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.43664e+32 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001101010100011010111000010111", b"00001101010100011010111000010111"), -- 0 + 6.46127e-31 = 6.46127e-31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01010110001100000101000111110101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.84665e+13 + inf = inf
	(b"10010000011010100100100011010100", b"00000000000000000000000000000000"),
	(b"11100011010010000001100101100010", b"11100011010010000001100101100010"), -- -4.62045e-29 + -3.69118e+21 = -3.69118e+21
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00111100001010101110010001011111", b"00000000000000000000000000000000"),
	(b"00000100010000000001100110010001", b"00111100001010101110010001011111"), -- 0.0104304 + 2.25812e-36 = 0.0104304
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101110100000011011001000110001", b"00101110100000011011001000110001"), -- 0 + 5.89789e-11 = 5.89789e-11
	(b"01001011000101111110010010101110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001011000101111110010010101110"), -- 9.95448e+06 + 0 = 9.95448e+06
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110100001100011011000111010001", b"01111111100000000000000000000000"), -- inf + 5.63137e+31 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111011111110001001011100111101", b"11111111100000000000000000000000"), -- -inf + -0.00758639 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000011011000000000010", b"10000000000000011011000000000010"), -- -0 + -1.54975e-40 = -1.54975e-40
	(b"01111101100110101010000101110001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.56924e+37 + inf = inf
	(b"10000000010010100110111011010001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000010010100110111011010001"), -- -6.83558e-39 + -0 = -6.83558e-39
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01101101100010101010010100011000", b"00000000000000000000000000000000"),
	(b"01000011010110001111011111100010", b"01101101100010101010010100011000"), -- 5.36356e+27 + 216.968 = 5.36356e+27
	(b"00010001100100000110011001001000", b"00000000000000000000000000000000"),
	(b"01110111000100001111001110010000", b"01110111000100001111001110010000"), -- 2.27822e-28 + 2.93996e+33 = 2.93996e+33
	(b"01000101010101010011100111100101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3411.62 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00100000011110101000111110001111", b"00000000000000000000000000000000"),
	(b"00100001001111011100011100101110", b"00100001011111000110101100010010"), -- 2.12233e-19 + 6.42993e-19 = 8.55226e-19
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10110000000000100110010110000000", b"00000000000000000000000000000000"),
	(b"11011010010100001010111000110011", b"11011010010100001010111000110011"), -- -4.7438e-10 + -1.46846e+16 = -1.46846e+16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110000101100010100010000110", b"00111110000101100010100010000110"), -- 0 + 0.146639 = 0.146639
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011111100111001001101110010000", b"01111111100000000000000000000000"), -- inf + 6.63259e-20 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00010001111110110111101101011001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.96768e-28 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00110110111111110111010101101101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00110110111111110111010101101101"), -- 7.61326e-06 + 0 = 7.61326e-06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10010001110011000011110111110110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.22237e-28 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010110101010010000110010111111", b"01111111100000000000000000000000"), -- inf + 9.29361e+13 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100011100001101100111110001101", b"01111111100000000000000000000000"), -- inf + 1.46162e-17 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11010100111110101001101100011011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11010100111110101001101100011011"), -- -8.61075e+12 + -0 = -8.61075e+12
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000011101010101101011100001011", b"11111111100000000000000000000000"), -- -inf + -341.68 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011001111100100010011101111010", b"11111111100000000000000000000000"), -- -inf + -2.50382e-23 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11011100110011111011000100011100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11011100110011111011000100011100"), -- -4.6768e+17 + -0 = -4.6768e+17
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000111111001", b"01111111100000000000000000000000"), -- inf + 7.07656e-43 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00111100110010111111001011101101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111100110010111111001011101101"), -- 0.0248961 + 0 = 0.0248961
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011110010000011110100011110011", b"11111111100000000000000000000000"), -- -inf + -1.02655e-20 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10101110011010010011110111011011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10101110011010010011110111011011"), -- -5.3033e-11 + -0 = -5.3033e-11
	(b"00000000000000000000000000001111", b"00000000000000000000000000000000"),
	(b"01111001110001100001011001100001", b"01111001110001100001011001100001"), -- 2.10195e-44 + 1.28566e+35 = 1.28566e+35
	(b"10001001111000000001101001011111", b"00000000000000000000000000000000"),
	(b"11110011111110011111110010001010", b"11110011111110011111110010001010"), -- -5.39508e-33 + -3.96119e+31 = -3.96119e+31
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110101000001100101110000101100", b"10110101000001100101110000101100"), -- -0 + -5.0053e-07 = -5.0053e-07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110111000101101101010000011100", b"00110111000101101101010000011100"), -- 0 + 8.99008e-06 = 8.99008e-06
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010000000010100101001100100110", b"11111111100000000000000000000000"), -- -inf + -9.28282e+09 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000010001000101000100011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000010001000101000100011"), -- 7.84238e-40 + 0 = 7.84238e-40
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000100100100011110010", b"01111111100000000000000000000000"), -- inf + 2.09839e-40 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111101010111100111110011010001", b"01111111100000000000000000000000"), -- inf + 1.84835e+37 = inf
	(b"00000000000000010111111111111111", b"00000000000000000000000000000000"),
	(b"01001011100010010010110101111001", b"01001011100010010010110101111001"), -- 1.37752e-40 + 1.79801e+07 = 1.79801e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011001010110010111111100000010", b"00011001010110010111111100000010"), -- 0 + 1.12443e-23 = 1.12443e-23
	(b"11101000100110010001100000001000", b"00000000000000000000000000000000"),
	(b"10111010000111001001111110000110", b"11101000100110010001100000001000"), -- -5.78372e+24 + -0.00059747 = -5.78372e+24
	(b"10011000000001111000011110000010", b"00000000000000000000000000000000"),
	(b"10101100100110110011111011100110", b"10101100100110110011111011100110"), -- -1.75168e-24 + -4.41235e-12 = -4.41235e-12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10101010100100000001110110110011", b"00000000000000000000000000000000"),
	(b"11010100000100111001111000100100", b"11010100000100111001111000100100"), -- -2.56001e-13 + -2.53605e+12 = -2.53605e+12
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000111001010000011101", b"10000000000000111001010000011101"), -- -0 + -3.2864e-40 = -3.2864e-40
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100111110010011101011000111001", b"11111111100000000000000000000000"), -- -inf + -1.90629e+24 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100101111010011010101010110100", b"11111111100000000000000000000000"), -- -inf + -1.37933e+23 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00001110101001001101110010011111", b"00000000000000000000000000000000"),
	(b"01001010011100100011101010000000", b"01001010011100100011101010000000"), -- 4.06416e-30 + 3.96867e+06 = 3.96867e+06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010000000000000010000001101001", b"11010000000000000010000001101001"), -- -0 + -8.59843e+09 = -8.59843e+09
	(b"01011110110111010101110001010011", b"00000000000000000000000000000000"),
	(b"01100001001000010010001100001110", b"01100001001010000000110111110001"), -- 7.97536e+18 + 1.85778e+20 = 1.93754e+20
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01010100001001000111001010100110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.82519e+12 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011110011110101100001000011100", b"00011110011110101100001000011100"), -- 0 + 1.3275e-20 = 1.3275e-20
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100110001100101101000011000100", b"10100110001100101101000011000100"), -- -0 + -6.20391e-16 = -6.20391e-16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10101100100010011001111101101011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.91147e-12 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110000110010000011100000100010", b"01111111100000000000000000000000"), -- inf + 1.45679e-09 = inf
	(b"10000000000000000000000000001100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000001100"), -- -1.68156e-44 + -0 = -1.68156e-44
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010001100101111100010110001111", b"01111111100000000000000000000000"), -- inf + 8.14818e+10 = inf
	(b"10100101101100100000001010110111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.08799e-16 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111101100010010100011100010011", b"11111101100010010100011100010011"), -- -0 + -2.28092e+37 = -2.28092e+37
	(b"00000000000000000011000111111011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.79296e-41 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010111111101001100100100110000", b"01010111111101001100100100110000"), -- 0 + 5.3829e+14 = 5.3829e+14
	(b"00100111100000110111111101000010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.64978e-15 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110010010101000101011101", b"01000000110010010101000101011101"), -- 0 + 6.29118 = 6.29118
	(b"10011000001000010110010010000101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10011000001000010110010010000101"), -- -2.08595e-24 + -0 = -2.08595e-24
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10101010110101011010100110001001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.7954e-13 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000001000001", b"01111111100000000000000000000000"), -- inf + 9.10844e-44 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100000011110111000101111011011", b"11111111100000000000000000000000"), -- -inf + -7.25033e+19 = -inf
	(b"01001101111010100100101101110001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001101111010100100101101110001"), -- 4.91352e+08 + 0 = 4.91352e+08
	(b"01001001001111011001111001100011", b"00000000000000000000000000000000"),
	(b"00101110100111001010011100111010", b"01001001001111011001111001100011"), -- 776678 + 7.12376e-11 = 776678
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011101001100111011101100100111", b"01011101001100111011101100100111"), -- 0 + 8.09437e+17 = 8.09437e+17
	(b"01011010001011111101100110010111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01011010001011111101100110010111"), -- 1.23743e+16 + 0 = 1.23743e+16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00100101001111101101011101110011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00100101001111101101011101110011"), -- 1.65529e-16 + 0 = 1.65529e-16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111001101110101001101000011011", b"01111111100000000000000000000000"), -- inf + 1.21112e+35 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101101100111100110100101101000", b"11101101100111100110100101101000"), -- -0 + -6.12826e+27 = -6.12826e+27
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01000011010011111101000101101001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000011010011111101000101101001"), -- 207.818 + 0 = 207.818
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01011011000011101000111010100111", b"00000000000000000000000000000000"),
	(b"00011001010011001001001111011111", b"01011011000011101000111010100111"), -- 4.01263e+16 + 1.05764e-23 = 4.01263e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100111101001111111000101101110", b"11111111100000000000000000000000"), -- -inf + -4.66136e-15 = -inf
	(b"10001100010101000010000110011010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.6342e-31 + -inf = -inf
	(b"11010100100001000101010011000001", b"00000000000000000000000000000000"),
	(b"11001001001111101111000111111001", b"11010100100001000101010011000010"), -- -4.54686e+12 + -782112 = -4.54686e+12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101011111111011010100101101011", b"11101011111111011010100101101011"), -- -0 + -6.13317e+26 = -6.13317e+26
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00011010000111000011111111000101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00011010000111000011111111000101"), -- 3.23116e-23 + 0 = 3.23116e-23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010011000001011001011010100100", b"00010011000001011001011010100100"), -- 0 + 1.68612e-27 = 1.68612e-27
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010011111000110000101101010001", b"11010011111000110000101101010001"), -- -0 + -1.95029e+12 = -1.95029e+12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11000010111101111010000110110100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000010111101111010000110110100"), -- -123.816 + -0 = -123.816
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101110100010001000100010100101", b"01111111100000000000000000000000"), -- inf + 6.20884e-11 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10111100010000111100110011110011", b"00000000000000000000000000000000"),
	(b"10101001111100101101001010110001", b"10111100010000111100110011110011"), -- -0.0119507 + -1.07835e-13 = -0.0119507
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101100000100011101100011010101", b"10101100000100011101100011010101"), -- -0 + -2.07261e-12 = -2.07261e-12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00010101111001011100010100000010", b"00000000000000000000000000000000"),
	(b"00110111100110110011110100001011", b"00110111100110110011110100001011"), -- 9.28032e-26 + 1.85059e-05 = 1.85059e-05
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000100010101010011111111110101", b"01000100010101010011111111110101"), -- 0 + 852.999 = 852.999
	(b"00000000000000000000000000010011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.66247e-44 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100101011001001010101001100100", b"01111111100000000000000000000000"), -- inf + 6.74902e+22 = inf
	(b"10100011100011000100110010011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100011100011000100110010011010"), -- -1.52113e-17 + -0 = -1.52113e-17
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011011100000011111100000110110", b"11111111100000000000000000000000"), -- -inf + -2.15017e-22 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000010100111110011111010110011", b"10000010100111110011111010110011"), -- -0 + -2.33989e-37 = -2.33989e-37
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01000000100001100100000101011001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.19548 + inf = inf
	(b"01011100101100001010010011100001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.97767e+17 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00011011101010000010100111100010", b"00000000000000000000000000000000"),
	(b"01001010010000000110101011010100", b"01001010010000000110101011010100"), -- 2.78203e-22 + 3.15256e+06 = 3.15256e+06
	(b"01000010101011100110001000001011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 87.1915 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11000100001000111011001100110010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -654.8 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101000100000101010110111011100", b"11111111100000000000000000000000"), -- -inf + -1.45083e-14 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010100000001000111110110101000", b"00010100000001000111110110101000"), -- 0 + 6.68908e-27 = 6.68908e-27
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010100100110111010011110111011", b"01010100100110111010011110111011"), -- 0 + 5.34827e+12 = 5.34827e+12
	(b"11111000001010100001101001111111", b"00000000000000000000000000000000"),
	(b"10101110011111101101000100100011", b"11111000001010100001101001111111"), -- -1.38004e+34 + -5.79387e-11 = -1.38004e+34
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000001111101100", b"00000000000000000000000000000000"),
	(b"00101010010110110111011111000100", b"00101010010110110111011111000100"), -- 1.4069e-42 + 1.94927e-13 = 1.94927e-13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10011001010100100111000101100010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10011001010100100111000101100010"), -- -1.08796e-23 + -0 = -1.08796e-23
	(b"10000001011000010100100101000011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.13785e-38 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00101000001001110111000101001111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.29493e-15 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00111110010000111110011101100100", b"00000000000000000000000000000000"),
	(b"00101000110010000011110010111010", b"00111110010000111110011101100100"), -- 0.191312 + 2.22308e-14 = 0.191312
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10110110111011101010010100001110", b"00000000000000000000000000000000"),
	(b"10011100101111011011000001110101", b"10110110111011101010010100001110"), -- -7.11217e-06 + -1.25526e-21 = -7.11217e-06
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000011010001100100001010100110", b"01111111100000000000000000000000"), -- inf + 5.82635e-37 = inf
	(b"10000000100001010001010001001001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000100001010001010001001001"), -- -1.22214e-38 + -0 = -1.22214e-38
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01000000100100000010001111101011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.50438 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100110111100111111101001110101", b"01100110111100111111101001110101"), -- 0 + 5.76078e+23 = 5.76078e+23
	(b"00000000000000000000000000000011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000011"), -- 4.2039e-45 + 0 = 4.2039e-45
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010011000011101011101010001000", b"01010011000011101011101010001000"), -- 0 + 6.13015e+11 = 6.13015e+11
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01011000011011011111011101111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000001000", b"01011000011011011111011101111011"), -- 1.04659e+15 + 1.12104e-44 = 1.04659e+15
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010100110000100010011011101111", b"10010100110000100010011011101111"), -- -0 + -1.96044e-26 = -1.96044e-26
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00010110100010100100111011010110", b"00000000000000000000000000000000"),
	(b"00000000000000000100101001101100", b"00010110100010100100111011010110"), -- 2.23449e-25 + 2.66975e-41 = 2.23449e-25
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01011000111111100100110000101110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.23683e+15 + inf = inf
	(b"01110111001111100110110111010000", b"00000000000000000000000000000000"),
	(b"01101001101010010111010111010101", b"01110111001111100110110111010000"), -- 3.86236e+33 + 2.56081e+25 = 3.86236e+33
	(b"00011110001110011001110100110111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.82633e-21 + inf = inf
	(b"10110000100010011000101011001100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110000100010011000101011001100"), -- -1.00075e-09 + -0 = -1.00075e-09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110011100011001001001111011010", b"01111111100000000000000000000000"), -- inf + 6.54615e-08 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011011010101001011100010010110", b"11011011010101001011100010010110"), -- -0 + -5.98756e+16 = -5.98756e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11100000000010100100000001100001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11100000000010100100000001100001"), -- -3.98483e+19 + -0 = -3.98483e+19
	(b"10011001011110000011010110011000", b"00000000000000000000000000000000"),
	(b"11001010100000111100011001010010", b"11001010100000111100011001010010"), -- -1.28321e-23 + -4.31799e+06 = -4.31799e+06
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01001011100011000110011000001000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001011100011000110011000001000"), -- 1.84023e+07 + 0 = 1.84023e+07
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000110110100010100101111001", b"00000000000000000000000000000000"),
	(b"01001010101000010110010011111011", b"01001010101000010110010011111011"), -- 2.0035e-38 + 5.28857e+06 = 5.28857e+06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000011000001000010100101011110", b"00000000000000000000000000000000"),
	(b"01111011000000100110000100000101", b"01111011000000100110000100000101"), -- 3.88388e-37 + 6.76966e+35 = 6.76966e+35
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011111001111011010011001001011", b"01111111100000000000000000000000"), -- inf + 4.01599e-20 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00101001000001111101111101010111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00101001000001111101111101010111"), -- 3.01697e-14 + 0 = 3.01697e-14
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111011011010101000100111001110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.21779e+36 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011111110010010111011111100101", b"01011111110010010111011111100101"), -- 0 + 2.90346e+19 = 2.90346e+19
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000001", b"01111111100000000000000000000000"), -- inf + 1.4013e-45 = inf
	(b"10100111001001100100110001000100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100111001001100100110001000100"), -- -2.30785e-15 + -0 = -2.30785e-15
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10001001010000000100111110101100", b"00000000000000000000000000000000"),
	(b"11110011110000000000011110100111", b"11110011110000000000011110100111"), -- -2.31486e-33 + -3.04284e+31 = -3.04284e+31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11101010110010010100011110101011", b"00000000000000000000000000000000"),
	(b"11100000000011001111110011101001", b"11101010110010010100011110101111"), -- -1.21666e+26 + -4.0637e+19 = -1.21666e+26
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10101011110111110100001110001011", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.58638e-12 + -inf = -inf
	(b"11010011100100011111110010000100", b"00000000000000000000000000000000"),
	(b"10011100100011101001101110010100", b"11010011100100011111110010000100"), -- -1.25401e+12 + -9.43699e-22 = -1.25401e+12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11101001110000011110101111100000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11101001110000011110101111100000"), -- -2.93046e+25 + -0 = -2.93046e+25
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000001110001110001010100101110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000001110001110001010100101110"), -- 7.31314e-38 + 0 = 7.31314e-38
	(b"01110100110011101001111011001011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.30961e+32 + inf = inf
	(b"10001010000110111011100001011001", b"00000000000000000000000000000000"),
	(b"10010000001011101101110100111110", b"10010000001011101110011011111010"), -- -7.49765e-33 + -3.44859e-29 = -3.44934e-29
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00100001010101100101001010011111", b"00000000000000000000000000000000"),
	(b"01100110000111100011001110110100", b"01100110000111100011001110110100"), -- 7.26154e-19 + 1.86772e+23 = 1.86772e+23
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100001001100010101010000010011", b"11111111100000000000000000000000"), -- -inf + -2.04446e+20 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110011101011100101101101001011", b"10110011101011100101101101001011"), -- -0 + -8.11911e-08 = -8.11911e-08
	(b"10111101001011000001110110100001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0.0420204 + -inf = -inf
	(b"00100000001001000111111011011001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.39333e-19 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11000011000110110001110000100000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -155.11 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10110011100010010001011110110101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.38387e-08 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100010011111101010110000010101", b"01111111100000000000000000000000"), -- inf + 1.17447e+21 = inf
	(b"00011101100000010110101100101110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.42568e-21 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10010101000010111000001110111101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.81747e-26 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011001000010011001111010000000", b"01011001000010011001111010000000"), -- 0 + 2.42102e+15 = 2.42102e+15
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10011010111011010100111110110110", b"00000000000000000000000000000000"),
	(b"11011011010011010101110001011010", b"11011011010011010101110001011010"), -- -9.81497e-23 + -5.78039e+16 = -5.78039e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11001000111000110100111001101101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001000111000110100111001101101"), -- -465523 + -0 = -465523
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11001111100001010101101110101111", b"00000000000000000000000000000000"),
	(b"10100000000111111111111110000010", b"11001111100001010101101110101111"), -- -4.47476e+09 + -1.35524e-19 = -4.47476e+09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010010100010101001110101101000", b"01111111100000000000000000000000"), -- inf + 2.97673e+11 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11100000000110101000010110000111", b"00000000000000000000000000000000"),
	(b"10111001010011000001101001011010", b"11100000000110101000010110000111"), -- -4.45378e+19 + -0.000194648 = -4.45378e+19
	(b"10111010110000101110011110110000", b"00000000000000000000000000000000"),
	(b"10011111101000111101110000000011", b"10111010110000101110011110110000"), -- -0.00148701 + -6.93972e-20 = -0.00148701
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010111010111110100010100111", b"11111111100000000000000000000000"), -- -inf + -3.32012e+16 = -inf
	(b"10101101000011011011100000110001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.05582e-12 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010000100111000111011001110011", b"11111111100000000000000000000000"), -- -inf + -6.17137e-29 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00010110010010100110011111100111", b"00000000000000000000000000000000"),
	(b"01111110010001001101101010100000", b"01111110010001001101101010100000"), -- 1.63502e-25 + 6.5416e+37 = 6.5416e+37
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111110111100001000010111101111", b"01111111100000000000000000000000"), -- inf + 1.59855e+38 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000010", b"11111111100000000000000000000000"), -- -inf + -2.8026e-45 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11101000010010000110010101001111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.78537e+24 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001010100110101011000000000010", b"01111111100000000000000000000000"), -- inf + 5.0688e+06 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000110000", b"00000000000000000000000000000000"),
	(b"10110110111010111010111011100111", b"10110110111010111010111011100111"), -- -6.72623e-44 + -7.02391e-06 = -7.02391e-06
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010100001011101100101011001110", b"11111111100000000000000000000000"), -- -inf + -8.82475e-27 = -inf
	(b"10000000000011000111101100010110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.14618e-39 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01010011100011000111110010000110", b"00000000000000000000000000000000"),
	(b"01011011111111000100101000011101", b"01011011111111000100101010101001"), -- 1.20677e+12 + 1.42026e+17 = 1.42028e+17
	(b"01010110111101101001100000110010", b"00000000000000000000000000000000"),
	(b"00011101010000100011000010111001", b"01010110111101101001100000110010"), -- 1.35567e+14 + 2.57009e-21 = 1.35567e+14
	(b"10000010011101000011011110001100", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.79422e-37 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001010010010011100110100000111", b"01111111100000000000000000000000"), -- inf + 3.30631e+06 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100010110001111101110000011111", b"11111111100000000000000000000000"), -- -inf + -5.41721e-18 = -inf
	(b"10010111110100111000001001100111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.36685e-24 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101110011100011001111111101100", b"01111111100000000000000000000000"), -- inf + 5.49391e-11 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111101100010000100001100101001", b"11111111100000000000000000000000"), -- -inf + -2.26405e+37 = -inf
	(b"10010011100000001111010011101000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.25532e-27 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011010001000011000110101001000", b"01111111100000000000000000000000"), -- inf + 3.34081e-23 = inf
	(b"10000111000000001100010101100010", b"00000000000000000000000000000000"),
	(b"11110101101110001100000101100100", b"11110101101110001100000101100100"), -- -9.68766e-35 + -4.68411e+32 = -4.68411e+32
	(b"10101111011010110000100000000010", b"00000000000000000000000000000000"),
	(b"11001000100011111011000110001000", b"11001000100011111011000110001000"), -- -2.1376e-10 + -294284 = -294284
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001010000101001001001100001110", b"01111111100000000000000000000000"), -- inf + 7.1536e-33 = inf
	(b"00111101110011101001100001000011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111101110011101001100001000011"), -- 0.100876 + 0 = 0.100876
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010010011010100101101110101", b"11011010010011010100101101110101"), -- -0 + -1.44463e+16 = -1.44463e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001010110111010111101111100100", b"11111111100000000000000000000000"), -- -inf + -7.25759e+06 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011110010110011001011001101110", b"11111111100000000000000000000000"), -- -inf + -1.1519e-20 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00100011001001101000001110101110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.02676e-18 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11110101100001000010000111101010", b"00000000000000000000000000000000"),
	(b"10011000001110011010100010111001", b"11110101100001000010000111101010"), -- -3.34996e+32 + -2.39959e-24 = -3.34996e+32
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11110011001001001000001000001001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110011001001001000001000001001"), -- -1.30337e+31 + -0 = -1.30337e+31
	(b"11001011000011110110100100111111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001011000011110110100100111111"), -- -9.39859e+06 + -0 = -9.39859e+06
	(b"10101010001001000101001100101110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10101010001001000101001100101110"), -- -1.4595e-13 + -0 = -1.4595e-13
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101001100000000110010011011001", b"01111111100000000000000000000000"), -- inf + 1.94023e+25 = inf
	(b"11110011011110101001111111101010", b"00000000000000000000000000000000"),
	(b"11101100110111100100100001010111", b"11110011011110101010011011011100"), -- -1.98565e+31 + -2.14979e+27 = -1.98587e+31
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100110100111010011111110000011", b"11111111100000000000000000000000"), -- -inf + -3.71292e+23 = -inf
	(b"00000000001110011101110011011111", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.31386e-39 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000010101000", b"00000000000000000000000010101000"), -- 0 + 2.35418e-43 = 2.35418e-43
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011111101001101100100111000011", b"01111111100000000000000000000000"), -- inf + 7.06375e-20 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000010", b"10000000000000000000000000000010"), -- -0 + -2.8026e-45 = -2.8026e-45
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110101101011100000111001101001", b"01111111100000000000000000000000"), -- inf + 4.41285e+32 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111010001010000111100100100011", b"10111010001010000111100100100011"), -- -0 + -0.000642674 = -0.000642674
	(b"00000001101100000000100000110011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.4664e-38 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111001000100101101011000001100", b"00000000000000000000000000000000"),
	(b"10101000010000010010110100101100", b"11111001000100101101011000001100"), -- -4.7651e+34 + -1.07234e-14 = -4.7651e+34
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11101011000001001011001010111001", b"00000000000000000000000000000000"),
	(b"10100001111101110010001101111000", b"11101011000001001011001010111001"), -- -1.60422e+26 + -1.67468e-18 = -1.60422e+26
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100101100011011001001010010101", b"01111111100000000000000000000000"), -- inf + 2.45589e-16 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01110110111100011000110000100111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01110110111100011000110000100111"), -- 2.44958e+33 + 0 = 2.44958e+33
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111011000000110011101101", b"01111111100000000000000000000000"), -- inf + 7.37658 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111101010011001101111100010000", b"11111111100000000000000000000000"), -- -inf + -1.702e+37 = -inf
	(b"01001011110110100111001110000101", b"00000000000000000000000000000000"),
	(b"00111100101110111011001011010101", b"01001011110110100111001110000101"), -- 2.86328e+07 + 0.0229124 = 2.86328e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101000000011110000101110000000", b"11111111100000000000000000000000"), -- -inf + -2.70204e+24 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000101101", b"11111111100000000000000000000000"), -- -inf + -6.30584e-44 = -inf
	(b"00001000110011111101101010110000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.25098e-33 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000011100010100000000000000101", b"01111111100000000000000000000000"), -- inf + 276 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001100110011110000111101111100", b"10001100110011110000111101111100"), -- -0 + -3.19027e-31 = -3.19027e-31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110101000011010010010110011101", b"10110101000011010010010110011101"), -- -0 + -5.25813e-07 = -5.25813e-07
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010101110101011110111010010110", b"00010101110101011110111010010110"), -- 0 + 8.64064e-26 = 8.64064e-26
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011011001000110110110101010110", b"11011011001000110110110101010110"), -- -0 + -4.60006e+16 = -4.60006e+16
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010110000111110101100110011", b"11011010110000111110101100110011"), -- -0 + -2.75731e+16 = -2.75731e+16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00101000010001000101100011101011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00101000010001000101100011101011"), -- 1.08995e-14 + 0 = 1.08995e-14
	(b"10001001101000111011011101001101", b"00000000000000000000000000000000"),
	(b"10111101110000101100011100100100", b"10111101110000101100011100100100"), -- -3.94132e-33 + -0.0951064 = -0.0951064
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001101100111110011100101100000", b"10001101100111110011100101100000"), -- -0 + -9.81294e-31 = -9.81294e-31
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00001000010001110111010100100100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00001000010001110111010100100100"), -- 6.00221e-34 + 0 = 6.00221e-34
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011101101110101001111101100000", b"01111111100000000000000000000000"), -- inf + 4.93986e-21 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100010100011100101101110", b"10111111100010100011100101101110"), -- -0 + -1.07988 = -1.07988
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001000011000100111101110011011", b"10001000011000100111101110011011"), -- -0 + -6.81547e-34 = -6.81547e-34
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01001010111001110111010011101001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000001", b"01001010111001110111010011101001"), -- 7.58437e+06 + 1.4013e-45 = 7.58437e+06
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111000110100001100011101110001", b"10111000110100001100011101110001"), -- -0 + -9.95536e-05 = -9.95536e-05
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110010100101100110000101110010", b"00110010100101100110000101110010"), -- 0 + 1.75066e-08 = 1.75066e-08
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00111000110011100001010001100100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111000110011100001010001100100"), -- 9.82664e-05 + 0 = 9.82664e-05
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101100101110101010100100111", b"00111101100101110101010100100111"), -- 0 + 0.0738929 = 0.0738929
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10001100000010100011010111010111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.06473e-31 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.00649e-45 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01100111000001001101001000111010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100111000001001101001000111010"), -- 6.2723e+23 + 0 = 6.2723e+23
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10100100100000011110011101111110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10100100100000011110011101111110"), -- -5.6337e-17 + -0 = -5.6337e-17
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101010010110100101001101010110", b"10101010010110100101001101010110"), -- -0 + -1.93912e-13 = -1.93912e-13
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101010110011110100110111101000", b"01111111100000000000000000000000"), -- inf + 3.68246e-13 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011000110000000000010110100010", b"01111111100000000000000000000000"), -- inf + 1.68904e+15 = inf
	(b"10110010011011000100000111010110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110010011011000100000111010110"), -- -1.3752e-08 + -0 = -1.3752e-08
	(b"11110011001000011100100000111001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110011001000011100100000111001"), -- -1.28177e+31 + -0 = -1.28177e+31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010101011000010111101110101111", b"01010101011000010111101110101111"), -- 0 + 1.54951e+13 = 1.54951e+13
	(b"11110111010000101011110000111010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110111010000101011110000111010"), -- -3.9497e+33 + -0 = -3.9497e+33
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010111010111111110101111000100", b"11010111010111111110101111000100"), -- -0 + -2.46204e+14 = -2.46204e+14
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001110111101111011000111011010", b"11001110111101111011000111011010"), -- -0 + -2.07781e+09 = -2.07781e+09
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100110110001111111100010100000", b"01111111100000000000000000000000"), -- inf + 1.38758e-15 = inf
	(b"01100100001001101010001001111010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100100001001101010001001111010"), -- 1.22955e+22 + 0 = 1.22955e+22
	(b"01010011101101100010100111001010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.56477e+12 + inf = inf
	(b"01111110101000000101101100110101", b"00000000000000000000000000000000"),
	(b"01101000100010000100000110101001", b"01111110101000000101101100110101"), -- 1.06575e+38 + 5.14762e+24 = 1.06575e+38
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001110100111010001011011010101", b"01111111100000000000000000000000"), -- inf + 1.31776e+09 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010010000100010010011100111000", b"00010010000100010010011100111000"), -- 0 + 4.58023e-28 = 4.58023e-28
	(b"10000000000000000000101110001000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000101110001000"), -- -4.13663e-42 + -0 = -4.13663e-42
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101101110011100111000000100", b"00111101101110011100111000000100"), -- 0 + 0.090725 = 0.090725
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111001010100100011111111100110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111001010100100011111111100110"), -- 6.82299e+34 + 0 = 6.82299e+34
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111001010111000111111101101110", b"00000000000000000000000000000000"),
	(b"10011010111111001010101111101100", b"11111001010111000111111101101110"), -- -7.15556e+34 + -1.04503e-22 = -7.15556e+34
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111001101111101011010111010011", b"10111001101111101011010111010011"), -- -0 + -0.000363751 = -0.000363751
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010100000010100111001101110001", b"01111111100000000000000000000000"), -- inf + 6.98999e-27 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010001011101010101110111100111", b"11010001011101010101110111100111"), -- -0 + -6.58652e+10 = -6.58652e+10
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000010001111101101111011110010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.4023e-37 + -inf = -inf
	(b"01000100011111100101110010000001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1017.45 + inf = inf
	(b"00010011011110011100101011010011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00010011011110011100101011010011"), -- 3.15282e-27 + 0 = 3.15282e-27
	(b"00000000000000011010000011101010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.49561e-40 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101111101111100010011111110011", b"00101111101111100010011111110011"), -- 0 + 3.45892e-10 = 3.45892e-10
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111011001111111011100111000110", b"11111111100000000000000000000000"), -- -inf + -9.95497e+35 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110001111001010101000011101001", b"11111111100000000000000000000000"), -- -inf + -2.27104e+30 = -inf
	(b"11010101110000001110011001110111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.6512e+13 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000111", b"11111111100000000000000000000000"), -- -inf + -9.80909e-45 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11100111101010111010010100110011", b"00000000000000000000000000000000"),
	(b"10111101011011000011011101100011", b"11100111101010111010010100110011"), -- -1.62114e+24 + -0.05767 = -1.62114e+24
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01100000110110111111110000010111", b"00000000000000000000000000000000"),
	(b"01111001101001110011110000000111", b"01111001101001110011110000000111"), -- 1.26813e+20 + 1.08541e+35 = 1.08541e+35
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111010101100001000111100001110", b"11111111100000000000000000000000"), -- -inf + -0.00134704 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100111101001010100001010001010", b"10100111101001010100001010001010"), -- -0 + -4.58688e-15 = -4.58688e-15
	(b"11111010011111000111111100100101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.27759e+35 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000110100010010000000010110000", b"11000110100010010000000010110000"), -- -0 + -17536.3 = -17536.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110010000111001100111100111100", b"01111111100000000000000000000000"), -- inf + 9.12751e-09 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001110100101000011101000101001", b"11111111100000000000000000000000"), -- -inf + -3.65408e-30 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101110101010011100111000101001", b"00101110101010011100111000101001"), -- 0 + 7.72185e-11 = 7.72185e-11
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000111111111111011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000111111111111011"), -- -4.59107e-41 + -0 = -4.59107e-41
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001000011010001111110000110", b"11111111100000000000000000000000"), -- -inf + -1.0663e+25 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000001111001100100001001010111", b"11111111100000000000000000000000"), -- -inf + -8.45838e-38 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011011111000011011100011101", b"01001011011111000011011100011101"), -- 0 + 1.65292e+07 = 1.65292e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001100100000100101001010111110", b"11111111100000000000000000000000"), -- -inf + -6.83269e+07 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00111101011110000001111100101011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0.0605766 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01000110100000001111001000111100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 16505.1 + inf = inf
	(b"01110011100110001011010110111111", b"00000000000000000000000000000000"),
	(b"00000100111001011100111011010010", b"01110011100110001011010110111111"), -- 2.41979e+31 + 5.40276e-36 = 2.41979e+31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101010010001001111010101011001", b"11101010010001001111010101011001"), -- -0 + -5.9527e+25 = -5.9527e+25
	(b"10001010001011100100100100000010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.39153e-33 + -inf = -inf
	(b"11011100011111001100010011010110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.84592e+17 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11010110000001011110011110001000", b"00000000000000000000000000000000"),
	(b"11101000101101000110111011000110", b"11101000101101000110111011000110"), -- -3.68074e+13 + -6.81656e+24 = -6.81656e+24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000011110011110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.73253e-42 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010101101100001011100110011101", b"11111111100000000000000000000000"), -- -inf + -7.13787e-26 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000101110101010010001001011000", b"11111111100000000000000000000000"), -- -inf + -6820.29 = -inf
	(b"10110101001000101100000111000010", b"00000000000000000000000000000000"),
	(b"11000010111011100011101011000011", b"11000010111011100011101011000011"), -- -6.06317e-07 + -119.115 = -119.115
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10101011100010010110010000001000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -9.7622e-13 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11100101011101001100101001011100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11100101011101001100101001011100"), -- -7.22494e+22 + -0 = -7.22494e+22
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01001100110000011101111011011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001100110000011101111011011010"), -- 1.01644e+08 + 0 = 1.01644e+08
	(b"11001001101010011001101010000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.38939e+06 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000001101010010111000110000011", b"11111111100000000000000000000000"), -- -inf + -6.22437e-38 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101111011001011011011100110000", b"11111111100000000000000000000000"), -- -inf + -2.08925e-10 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101000011011100100011001010001", b"01111111100000000000000000000000"), -- inf + 4.50088e+24 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01110110101001100110011001010101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.68749e+33 + inf = inf
	(b"01000011111100101110111111101110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 485.874 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01100001100011011101011100111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100001100011011101011100111011"), -- 3.27062e+20 + 0 = 3.27062e+20
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011110010110011101011110110111", b"01011110010110011101011110110111"), -- 0 + 3.9243e+18 = 3.9243e+18
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000001000000", b"01111111100000000000000000000000"), -- inf + 8.96831e-44 = inf
	(b"00111001111110101100000101101001", b"00000000000000000000000000000000"),
	(b"00000000001101000000010110100011", b"00111001111110101100000101101001"), -- 0.000478278 + 4.77747e-39 = 0.000478278
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11110000001111110010100010111110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110000001111110010100010111110"), -- -2.36644e+29 + -0 = -2.36644e+29
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01100001011100101011110110110001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100001011100101011110110110001"), -- 2.79861e+20 + 0 = 2.79861e+20
	(b"10011001000000000101001000010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.63402e-24 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111011001000001011110000110010", b"01111111100000000000000000000000"), -- inf + 8.34585e+35 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001101001001100101110011000011", b"01001101001001100101110011000011"), -- 0 + 1.74444e+08 = 1.74444e+08
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001111101101110001001000001111", b"11111111100000000000000000000000"), -- -inf + -1.80521e-29 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01100100001011100101011100010001", b"00000000000000000000000000000000"),
	(b"00111100001010100011101011101111", b"01100100001011100101011100010001"), -- 1.2864e+22 + 0.01039 = 1.2864e+22
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011111001000111100100110101111", b"11011111001000111100100110101111"), -- -0 + -1.18022e+19 = -1.18022e+19
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011000111111101111111", b"01111111100000000000000000000000"), -- inf + 3.69528 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01100111011000111101001010000101", b"00000000000000000000000000000000"),
	(b"00001111100110110001001110000110", b"01100111011000111101001010000101"), -- 1.07586e+24 + 1.52917e-29 = 1.07586e+24
	(b"10000101100010000101011001001111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000101100010000101011001001111"), -- -1.28211e-35 + -0 = -1.28211e-35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111011001000100110100111110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -3.03465e+38 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000101110111011100100000111010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000101110111011100100000111010"), -- -2.08563e-35 + -0 = -2.08563e-35
	(b"00010100111100000001011010001110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.42427e-26 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01011111101101100011001011110100", b"01111111100000000000000000000000"), -- inf + 2.62576e+19 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001001010001001111001000010011", b"01111111100000000000000000000000"), -- inf + 806689 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00100011111010110001101110001100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.54904e-17 + inf = inf
	(b"10111011100011100101111010101011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111011100011100101111010101011"), -- -0.00434478 + -0 = -0.00434478
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001101101110110110000000100010", b"11111111100000000000000000000000"), -- -inf + -3.92955e+08 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100110110111011000011001111111", b"11100110110111011000011001111111"), -- -0 + -5.23062e+23 = -5.23062e+23
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10011110011000000001010000101010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.18626e-20 + -inf = -inf
	(b"11111101101001011000001111100011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111101101001011000001111100011"), -- -2.75009e+37 + -0 = -2.75009e+37
	(b"01011110011101110100110100101000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.45499e+18 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11110000011111000110001111100111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110000011111000110001111100111"), -- -3.12444e+29 + -0 = -3.12444e+29
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10111100100010101111101100010101", b"00000000000000000000000000000000"),
	(b"11110000110000110011001011010001", b"11110000110000110011001011010001"), -- -0.0169654 + -4.83288e+29 = -4.83288e+29
	(b"10010001010111001100111111001000", b"00000000000000000000000000000000"),
	(b"10101101000100100101000100001111", b"10101101000100100101000100001111"), -- -1.7419e-28 + -8.31714e-12 = -8.31714e-12
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000110101101001100001101010011", b"00000000000000000000000000000000"),
	(b"10111011111000011010011100000101", b"10111011111000011010011100000101"), -- -6.79955e-35 + -0.00688637 = -0.00688637
	(b"11010000001011101100011100100101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.17291e+10 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010000000101001110011110000101", b"01111111100000000000000000000000"), -- inf + 2.93662e-29 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001101001000110011000110110000", b"01111111100000000000000000000000"), -- inf + 1.71121e+08 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010001010100111011001011110", b"11011010001010100111011001011110"), -- -0 + -1.19952e+16 = -1.19952e+16
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001110111001110110100110110101", b"01111111100000000000000000000000"), -- inf + 5.70477e-30 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010110110001000111101101110111", b"01111111100000000000000000000000"), -- inf + 3.17434e-25 = inf
	(b"00110111010001000010001000000100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00110111010001000010001000000100"), -- 1.16904e-05 + 0 = 1.16904e-05
	(b"11100101110000000100100100001100", b"00000000000000000000000000000000"),
	(b"10101001000110110000000010101000", b"11100101110000000100100100001100"), -- -1.13505e+23 + -3.44175e-14 = -1.13505e+23
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10011011100111011101001001001110", b"00000000000000000000000000000000"),
	(b"10010111101010000111001100110000", b"10011011100111100111101011000001"), -- -2.61094e-22 + -1.08858e-24 = -2.62182e-22
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10001000001101000100110110110110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.42581e-34 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011101011011100101110000111100", b"10011101011011100101110000111100"), -- -0 + -3.15467e-21 = -3.15467e-21
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00101000001100000010000001111001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.777e-15 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11011010001000001000011010000001", b"11011010001000001000011010000001"), -- -0 + -1.1296e+16 = -1.1296e+16
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01101000010010110000100101011101", b"01101000010010110000100101011101"), -- 0 + 3.83525e+24 = 3.83525e+24
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110110100100101000011111111101", b"11111111100000000000000000000000"), -- -inf + -4.36697e-06 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000011010010", b"00000000000000000000000000000000"),
	(b"00101011010100010111110010010001", b"00101011010100010111110010010001"), -- 2.94273e-43 + 7.44246e-13 = 7.44246e-13
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01011110110101000011101110001011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 7.64648e+18 + inf = inf
	(b"01100110001010000001100011010111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100110001010000001100011010111"), -- 1.98454e+23 + 0 = 1.98454e+23
	(b"00101101001110001000101100010100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.04901e-11 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01101010000011000110110110101010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101010000011000110110110101010"), -- 4.24419e+25 + 0 = 4.24419e+25
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101110011001111000001111", b"01111111100000000000000000000000"), -- inf + 92.8087 = inf
	(b"10011110010000001000000011110100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10011110010000001000000011110100"), -- -1.01911e-20 + -0 = -1.01911e-20
	(b"11010101111100100101000111010110", b"00000000000000000000000000000000"),
	(b"11000100100001100010101110101001", b"11010101111100100101000111010110"), -- -3.33042e+13 + -1073.36 = -3.33042e+13
	(b"11101010001000100100010110101000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11101010001000100100010110101000"), -- -4.90437e+25 + -0 = -4.90437e+25
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11011101010111001100111010111000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11011101010111001100111010111000"), -- -9.94429e+17 + -0 = -9.94429e+17
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001101111101100000110101110101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001101111101100000110101110101"), -- -5.1601e+08 + -0 = -5.1601e+08
	(b"01111010110001000111100100101110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111010110001000111100100101110"), -- 5.10074e+35 + 0 = 5.10074e+35
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00100001001000110010001110111101", b"00100001001000110010001110111101"), -- 0 + 5.52738e-19 = 5.52738e-19
	(b"00000000010000000101011001010011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000010000000101011001010011"), -- 5.90844e-39 + 0 = 5.90844e-39
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001101001111101010110010011100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001101001111101010110010011100"), -- 1.99936e+08 + 0 = 1.99936e+08
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01100010010111110011010100110001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01100010010111110011010100110001"), -- 1.02936e+21 + 0 = 1.02936e+21
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101100100001001000100101110100", b"10101100100001001000100101110100"), -- -0 + -3.76693e-12 = -3.76693e-12
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100100011011000111000000111010", b"11111111100000000000000000000000"), -- -inf + -5.12694e-17 = -inf
	(b"00110100001101111000100111111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00110100001101111000100111111011"), -- 1.70934e-07 + 0 = 1.70934e-07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00011111101110101110000010010011", b"00000000000000000000000000000000"),
	(b"00110001011101100010100000011001", b"00110001011101100010100000011001"), -- 7.91456e-20 + 3.58205e-09 = 3.58205e-09
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001100110011111111011111", b"11111111100000000000000000000000"), -- -inf + -4.70652e-39 = -inf
	(b"11110001110001111011101100011101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.97804e+30 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"00111111110010000000000100111101", b"00000000000000000000000000000000"),
	(b"01101011001100100111011011001110", b"01101011001100100111011011001110"), -- 1.56254 + 2.1575e+26 = 2.1575e+26
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010101011011110001101001111001", b"00010101011011110001101001111001"), -- 0 + 4.82865e-26 = 4.82865e-26
	(b"11101100100110010111010000111101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11101100100110010111010000111101"), -- -1.48412e+27 + -0 = -1.48412e+27
	(b"11110000010000100111100100110000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110000010000100111100100110000"), -- -2.40746e+29 + -0 = -2.40746e+29
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10110101001000000010100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110101001000000010100110011010"), -- -5.96652e-07 + -0 = -5.96652e-07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11110011000110011111011111000000", b"11111111100000000000000000000000"), -- -inf + -1.21986e+31 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.4013e-45 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100011100011111000011111001101", b"10100011100011111000011111001101"), -- -0 + -1.55616e-17 = -1.55616e-17
	(b"11011100111010111011111110001011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11011100111010111011111110001011"), -- -5.30858e+17 + -0 = -5.30858e+17
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11100101111010001101101111011101", b"11111111100000000000000000000000"), -- -inf + -1.37456e+23 = -inf
	(b"10001110100111110010001111001110", b"00000000000000000000000000000000"),
	(b"10000000000000000000100010000010", b"10001110100111110010001111001110"), -- -3.9231e-30 + -3.05203e-42 = -3.9231e-30
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001001111001010111010010111011", b"00001001111001010111010010111011"), -- 0 + 5.52395e-33 = 5.52395e-33
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000001011010101011010001100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.16364e-39 + inf = inf
	(b"10111101001010001110111110000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0.041244 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100100001110110110110100001101", b"11111111100000000000000000000000"), -- -inf + -4.06415e-17 = -inf
	(b"01111001000100111001111111101010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 4.79069e+34 + inf = inf
	(b"10001110110100010001010110111011", b"00000000000000000000000000000000"),
	(b"10110010000100010100001110100111", b"10110010000100010100001110100111"), -- -5.15434e-30 + -8.45549e-09 = -8.45549e-09
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10010010111001111010110111111111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.4621e-27 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000111010", b"11111111100000000000000000000000"), -- -inf + -8.12753e-44 = -inf
	(b"00100000011010101100101110011101", b"00000000000000000000000000000000"),
	(b"00001000000011101110101100011000", b"00100000011010101100101110011101"), -- 1.98879e-19 + 4.30079e-34 = 1.98879e-19
	(b"11000111000011010010011000001000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -36134 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101100000111000011101100110010", b"00101100000111000011101100110010"), -- 0 + 2.22018e-12 = 2.22018e-12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111110111101001000001010101001", b"11111110111101001000001010101001"), -- -0 + -1.62505e+38 = -1.62505e+38
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101011010111111000010110011110", b"10101011010111111000010110011110"), -- -0 + -7.94109e-13 = -7.94109e-13
	(b"10011000111100101001011101100000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -6.27084e-24 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001111101101011111100011111011", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 6.10599e+09 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111000111000001000000111110011", b"11111000111000001000000111110011"), -- -0 + -3.64284e+34 = -3.64284e+34
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101101111010011110011100010011", b"10101101111010011110011100010011"), -- -0 + -2.65917e-11 = -2.65917e-11
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00010111101011100101111100011111", b"00010111101011100101111100011111"), -- 0 + 1.12685e-24 = 1.12685e-24
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01000100011001000001111010100110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 912.479 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01001100000100011001101110000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001100000100011001101110000000"), -- 3.81701e+07 + 0 = 3.81701e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000001011011000110100001100", b"10000000001011011000110100001100"), -- -0 + -4.1832e-39 = -4.1832e-39
	(b"11111101100100101001110010001001", b"00000000000000000000000000000000"),
	(b"10110100100000010011101001001111", b"11111101100100101001110010001001"), -- -2.436e+37 + -2.40705e-07 = -2.436e+37
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01000000101010111101010111011100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000000101010111101010111011100"), -- 5.36986 + 0 = 5.36986
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101111011001000010100110101100", b"11111111100000000000000000000000"), -- -inf + -2.07513e-10 = -inf
	(b"10110001000110011110001000011000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10110001000110011110001000011000"), -- -2.23929e-09 + -0 = -2.23929e-09
	(b"10000000000000000000000000000001", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.4013e-45 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001110010111011111111011000000", b"00001110010111011111111011000000"), -- 0 + 2.7363e-30 = 2.7363e-30
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10010111000100110000111110000010", b"11111111100000000000000000000000"), -- -inf + -4.75178e-25 = -inf
	(b"00110001110110001101101010010001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00110001110110001101101010010001"), -- 6.31128e-09 + 0 = 6.31128e-09
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100111010110000100110111100111", b"01100111010110000100110111100111"), -- 0 + 1.02147e+24 = 1.02147e+24
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001101001101000011000100111", b"11101001101001101000011000100111"), -- -0 + -2.51644e+25 = -2.51644e+25
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000001", b"01111111100000000000000000000000"), -- inf + 1.4013e-45 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000001", b"00000000000000000000000000000001"), -- 0 + 1.4013e-45 = 1.4013e-45
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000111101110001100100010", b"00000000000000000000000000000000"),
	(b"10011011010111001000111100111101", b"10011011010111001000111100111101"), -- -2.83654e-39 + -1.82443e-22 = -1.82443e-22
	(b"00110100000111110111010101101101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.48507e-07 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00100111100111001010101110100000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00100111100111001010101110100000"), -- 4.34848e-15 + 0 = 4.34848e-15
	(b"00100100000011000010000010011001", b"00000000000000000000000000000000"),
	(b"00010011000001111000011111011111", b"00100100000011000010000010011001"), -- 3.03853e-17 + 1.71064e-27 = 3.03853e-17
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110111011111111000110111111001", b"00110111011111111000110111111001"), -- 0 + 1.52322e-05 = 1.52322e-05
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111011100000011100000010010011", b"01111111100000000000000000000000"), -- inf + 0.00395972 = inf
	(b"00100000101000000001110010101110", b"00000000000000000000000000000000"),
	(b"00011110010000000111101101010000", b"00100000101001100010000010001000"), -- 2.7124e-19 + 1.01899e-20 = 2.8143e-19
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01110010110101000000001011001010", b"01110010110101000000001011001010"), -- 0 + 8.39862e+30 = 8.39862e+30
	(b"01101101100010110000011101000001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101101100010110000011101000001"), -- 5.3784e+27 + 0 = 5.3784e+27
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00011111110001001001000101100100", b"01111111100000000000000000000000"), -- inf + 8.32498e-20 = inf
	(b"11110011011111111001011111011001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11110011011111111001011111011001"), -- -2.02502e+31 + -0 = -2.02502e+31
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111100000000101100010001100010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.71593e+36 + inf = inf
	(b"01111110000101010001000100010011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111110000101010001000100010011"), -- 4.95359e+37 + 0 = 4.95359e+37
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111010011110010011011011100100", b"11111010011110010011011011100100"), -- -0 + -3.23499e+35 = -3.23499e+35
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111010010110011110100101100010", b"01111010010110011110100101100010"), -- 0 + 2.82865e+35 = 2.82865e+35
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01100011000110101011111001000101", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.85451e+21 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101001011110001101001100011111", b"11111111100000000000000000000000"), -- -inf + -1.88007e+25 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01100100100011001000110111001001", b"01111111100000000000000000000000"), -- inf + 2.07421e+22 = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10001001101001010001010010100101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10001001101001010001010010100101"), -- -3.97417e-33 + -0 = -3.97417e-33
	(b"01001010100001110000011101101100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001010100001110000011101101100"), -- 4.42463e+06 + 0 = 4.42463e+06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10010101010001010001100010110000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10010101010001010001100010110000"), -- -3.98033e-26 + -0 = -3.98033e-26
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"00000000000001101111101010010111", b"00000000000000000000000000000000"),
	(b"01101110100111111101010011000000", b"01101110100111111101010011000000"), -- 6.40908e-40 + 2.47327e+28 = 2.47327e+28
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001110001100010000011111001100", b"10001110001100010000011111001100"), -- -0 + -2.18207e-30 = -2.18207e-30
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"11100100010100001101101000100011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11100100010100001101101000100011"), -- -1.54106e+22 + -0 = -1.54106e+22
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10100001100011100100110110110101", b"10100001100011100100110110110101"), -- -0 + -9.64286e-19 = -9.64286e-19
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00001000000000001000011110111010", b"01111111100000000000000000000000"), -- inf + 3.86781e-34 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10101000100011101000001101101100", b"00000000000000000000000000000000"),
	(b"10100111001101010010011101001001", b"10101000101001010010100001010101"), -- -1.58222e-14 + -2.51401e-15 = -1.83362e-14
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010101110111101111001110010111", b"11111111100000000000000000000000"), -- -inf + -3.06422e+13 = -inf
	(b"10011011000110110110100100010110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10011011000110110110100100010110"), -- -1.28553e-22 + -0 = -1.28553e-22
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000010010101100100010111100111", b"00000010010101100100010111100111"), -- 0 + 1.57423e-37 = 1.57423e-37
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000001", b"00000000000000000000000000000001"), -- 0 + 1.4013e-45 = 1.4013e-45
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010011000010101011000101110110", b"11111111100000000000000000000000"), -- -inf + -5.95683e+11 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10011000101000110100100011101111", b"11111111100000000000000000000000"), -- -inf + -4.22082e-24 = -inf
	(b"01110010111010110010010111010111", b"00000000000000000000000000000000"),
	(b"00101010101001100011100001011100", b"01110010111010110010010111010111"), -- 9.31516e+30 + 2.95266e-13 = 9.31516e+30
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10101000110111010111000100101110", b"10101000110111010111000100101110"), -- -0 + -2.4585e-14 = -2.4585e-14
	(b"10011000100010110010111000001111", b"00000000000000000000000000000000"),
	(b"10010101110100101101111111000111", b"10011000100011100111100110001110"), -- -3.59772e-24 + -8.51714e-26 = -3.68289e-24
	(b"00101010110010110110001100101100", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 3.61289e-13 + inf = inf
	(b"10000000000000000000011110001010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.70451e-42 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11111000010010011010011110101000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -1.63602e+34 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01010011100001011101001011011100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01010011100001011101001011011100"), -- 1.14954e+12 + 0 = 1.14954e+12
	(b"00111001011100110110001100010001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111001011100110110001100010001"), -- 0.000232112 + 0 = 0.000232112
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111110100000010100100010111101", b"01111111100000000000000000000000"), -- inf + 8.5924e+37 = inf
	(b"01011001011011110001000001110011", b"00000000000000000000000000000000"),
	(b"00011111111001000001000000010100", b"01011001011011110001000001110011"), -- 4.20566e+15 + 9.65884e-20 = 4.20566e+15
	(b"11100110110001000101011010100111", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -4.63591e+23 + -inf = -inf
	(b"00001110000001010101111101111000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.64395e-30 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00101100011010011100001111010011", b"01111111100000000000000000000000"), -- inf + 3.322e-12 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111010111111110101101010010001", b"11111010111111110101101010010001"), -- -0 + -6.62936e+35 = -6.62936e+35
	(b"10001101010100100110010101110111", b"00000000000000000000000000000000"),
	(b"10111000010001110000101010011111", b"10111000010001110000101010011111"), -- -6.48334e-31 + -4.74552e-05 = -4.74552e-05
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"11100100100110010100000001000101", b"00000000000000000000000000000000"),
	(b"11110110010111110011101011011101", b"11110110010111110011101011011101"), -- -2.26159e+22 + -1.13191e+33 = -1.13191e+33
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01000001111011000001100110101010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000001111011000001100110101010"), -- 29.5125 + 0 = 29.5125
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11001011111100111000111110100000", b"00000000000000000000000000000000"),
	(b"10001111010100000110111000010100", b"11001011111100111000111110100000"), -- -3.1924e+07 + -1.02764e-29 = -3.1924e+07
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"01000010101000101011011110110000", b"00000000000000000000000000000000"),
	(b"00111011100000101111100110111100", b"01000010101000101011100110111100"), -- 81.3588 + 0.00399706 = 81.3628
	(b"11111100011111111110011010010101", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -5.31485e+36 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10110100010011000101100111010011", b"10110100010011000101100111010011"), -- -0 + -1.90317e-07 = -1.90317e-07
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111101010101100000001000011111", b"01111111100000000000000000000000"), -- inf + 1.77791e+37 = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00111000110101100001001001100010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0.000102077 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10111010000111000000001011011101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111010000111000000001011011101"), -- -0.000595135 + -0 = -0.000595135
	(b"11000011000100011100010001011010", b"00000000000000000000000000000000"),
	(b"11100101111110100011010101010010", b"11100101111110100011010101010010"), -- -145.767 + -1.47697e+23 = -1.47697e+23
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00100001101000111001001110101011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00100001101000111001001110101011"), -- 1.10844e-18 + 0 = 1.10844e-18
	(b"11101010110111101101101110011000", b"00000000000000000000000000000000"),
	(b"10010000001100101100110001001111", b"11101010110111101101101110011000"), -- -1.34709e+26 + -3.52617e-29 = -1.34709e+26
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00000000000000100000100010010110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.86751e-40 + inf = inf
	(b"01111100111010111011101101101000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 9.79193e+36 + inf = inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111000010100011110010110000100", b"00111000010100011110010110000100"), -- 0 + 5.00432e-05 = 5.00432e-05
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111010010011110001100100110000", b"11111010010011110001100100110000"), -- -0 + -2.68829e+35 = -2.68829e+35
	(b"00110001000101100100011111111110", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 2.18688e-09 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -0 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- inf + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000010110011", b"00000000000000000000000000000000"),
	(b"10011010111011011011101001101001", b"10011010111011011011101001101001"), -- -2.50832e-43 + -9.83221e-23 = -9.83221e-23
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111100101110001001101010010010", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -7.66814e+36 + -inf = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11010010100001011101101110010110", b"11010010100001011101101110010110"), -- -0 + -2.87457e+11 = -2.87457e+11
	(b"01101011111000001011011100110010", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.43329e+26 + inf = inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111010100010110001101010001000", b"11111111100000000000000000000000"), -- -inf + -0.00106128 = -inf
	(b"11111010000111111000010101110001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11111010000111111000010101110001"), -- -2.0707e+35 + -0 = -2.0707e+35
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10001111010110000001011110011111", b"10001111010110000001011110011111"), -- -0 + -1.06542e-29 = -1.06542e-29
	(b"01101110010100011100101000111001", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 1.62317e+28 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01111111100000000000000000000000"), -- inf + 0 = inf
	(b"10110010110100011101101101011000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -2.44305e-08 + -inf = -inf
	(b"00010000100000011111110100010000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 5.12714e-29 + inf = inf
	(b"01111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01010011101000010100011011001111", b"01111111100000000000000000000000"), -- inf + 1.38536e+12 = inf
	(b"01010010001001001010100110000111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01010010001001001010100110000111"), -- 1.76805e+11 + 0 = 1.76805e+11
	(b"10101101000101101111111011111110", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -8.58313e-12 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"00011100100000011110100000000000", b"00000000000000000000000000000000"),
	(b"01001101101000011000000011001111", b"01001101101000011000000011001111"), -- 8.59647e-22 + 3.38697e+08 = 3.38697e+08
	(b"10000110110001011101110001100111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000110110001011101110001100111"), -- -7.4427e-35 + -0 = -7.4427e-35
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11101000100101011100011011000010", b"11111111100000000000000000000000"), -- -inf + -5.65839e+24 = -inf
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00110011000101100011010011011000", b"00110011000101100011010011011000"), -- 0 + 3.49727e-08 = 3.49727e-08
	(b"01101101100011001110010010101100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01101101100011001110010010101100"), -- 5.45054e+27 + 0 = 5.45054e+27
	(b"11111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -inf + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11111111100000000000000000000000", b"11111111100000000000000000000000"), -- -0 + -inf = -inf
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01111111100000000000000000000000", b"01111111100000000000000000000000"), -- 0 + inf = inf

	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000111000101110110101000011111", b"11001011101000111000101101010101"), -- -2.14748e+07 + 38762.1 = -2.14361e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001000001101000011000001011111", b"00000000000000000000000000000000"),
	(b"01000111000001011110011101010100", b"01001000010101011010101000110100"), -- 184513 + 34279.3 = 218793
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111101110011001100110011010", b"11001011101000111101011100001001"), -- -2.14748e+07 + 1.45 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11000010100001000101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011011101001"), -- -66.17 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001000111100100001110011011010", b"11001000111100100001110011011010"), -- -0 + -495847 = -495847
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111110100110011001100110011010"), -- -0.3 + -0 = -0.3
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0.01 = 2.14748e+07
	(b"01000111111110000100001111101111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000111111110000100001111101111"), -- 127112 + 0 = 127112
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001010101100101011110000000101", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011011011100101000000010010"), -- 5.85677e+06 + -2.14748e+07 = -1.56181e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11000011100011100111110101110001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000011100011100111110101110001"), -- -284.98 + -0 = -284.98
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0.47 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"00111110010000101000111101011100"), -- 0 + 0.19 = 0.19
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0.03 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0.15 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11000010101111011000111101011100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000010101111011000111101011100"), -- -94.78 + -0 = -94.78
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011000100010101000110000111", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001011000100010101000110000111"), -- -9.52359e+06 + -0 = -9.52359e+06
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001000001010000001010001110010", b"11001000001010000001010001110010"), -- -0 + -172114 = -172114
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001000110010001111011000110011", b"01001011101000001011001100110001"), -- 2.14748e+07 + -411570 = 2.10633e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01000000101100100011110101110001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000000101100100011110101110001"), -- 5.57 + 0 = 5.57
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000101101011000000111111010111", b"01000101101011000000111111010111"), -- 0 + 5505.98 = 5505.98
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011011010111011000100010001", b"11001011011010111011000100010001"), -- -0 + -1.54463e+07 = -1.54463e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100101000111101011100", b"01000000011100101000111101011100"), -- 0 + 3.79 = 3.79
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001010001001011011011010011010", b"01001010001001011011011010011010"), -- 0 + 2.71505e+06 = 2.71505e+06
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000010001101000100011110101110", b"01001011101000111101011011110011"), -- 2.14748e+07 + -45.07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11000011000101000101010001111011", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011011000000"), -- -148.33 + 2.14748e+07 = 2.14747e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000111100110001000110100000011", b"01001011101000110011111001111101"), -- 2.14748e+07 + -78106 = 2.13967e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000011010011100101011100001010", b"01001011101000111101011010100011"), -- 2.14748e+07 + -206.34 = 2.14746e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"10111101011101011100001010001111"), -- -0 + -0.06 = -0.06
	(b"11000110001111000110001001001000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111011111101111110"), -- -12056.6 + 2.14748e+07 = 2.14628e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001010011100000011000100110111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01001010011100000011000100110111"), -- 3.93531e+06 + 0 = 3.93531e+06
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01000111011001101011000000101001", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000110110001110110010"), -- 59056.2 + -2.14748e+07 = -2.14158e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001001001111110011111111001010", b"11001011100111011101110100001100"), -- -2.14748e+07 + 783357 = -2.06915e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111010111101011100001010010"), -- -0 + -0.87 = -0.87
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01000011010001101001111010111000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000011010001101001111010111000"), -- 198.62 + 0 = 198.62
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111101111101011100001010001111"), -- 0.12 + 0 = 0.12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000111100110010011011010011100", b"11000111100110010011011010011100"), -- -0 + -78445.2 = -78445.2
	(b"11001000101100110100100010000101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001000101100110100100010000101"), -- -367172 + -0 = -367172
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01000010101100110111000010100100", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011011011101"), -- 89.72 + -2.14748e+07 = -2.14747e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001001100001101100101001101100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001001100001101100101001101100"), -- -1.10421e+06 + -0 = -1.10421e+06
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000100110000100100100111101100", b"11000100110000100100100111101100"), -- -0 + -1554.31 = -1554.31
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001001000100110111100100010011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11001001000100110111100100010011"), -- -604049 + -0 = -604049
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001001100100011110001000001011", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011100110101011100011101001"), -- 1.19507e+06 + -2.14748e+07 = -2.02798e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11000101001111110000110011110110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000101001111110000110011110110"), -- -3056.81 + -0 = -3056.81
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0.59 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11000001110100000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000001110100000000000000000000"), -- -26 + -0 = -26
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000100010101101000110000101001", b"01000100010101101000110000101001"), -- 0 + 858.19 = 858.19
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001000000000100100000100010010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000101101001010001000"), -- -133380 + 2.14748e+07 = 2.13415e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111101100011110101110000101001"), -- -0.07 + -0 = -0.07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11000001100001010101110000101001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000001100001010101110000101001"), -- -16.67 + -0 = -16.67
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000111100101011000010000011100", b"01000111100101011000010000011100"), -- 0 + 76552.2 = 76552.2
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001001001011101110101100010110", b"11001001001011101110101100010110"), -- -0 + -716465 = -716465
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000100110001000011111100001010", b"11001011101000111101001111111001"), -- -2.14748e+07 + 1569.97 = -2.14733e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101011100110011001100110", b"11000000101011100110011001100110"), -- -0 + -5.45 = -5.45
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000110100000001100100011001101", b"01000110100000001100100011001101"), -- 0 + 16484.4 = 16484.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11000000100101110000101000111101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000100101110000101000111101"), -- -4.72 + -0 = -4.72
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000001111110101100110011001101", b"01001011101000111101011011111010"), -- 2.14748e+07 + -31.35 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110111000010100011110101110", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0.44 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111000101000111101011100001"), -- 0 + 0.58 = 0.58
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01000101001111110001110001111011", b"00000000000000000000000000000000"),
	(b"01000011000000001111100001010010", b"01000101010001110010110000000000"), -- 3057.78 + 128.97 = 3186.75
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001000101101000101111001010111", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000010000010110010001"), -- -369395 + 2.14748e+07 = 2.11054e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111111001010111000010100011111"), -- 0.67 + 0 = 0.67
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001010011100100010100011100001", b"01001011100001011001000111101110"), -- 2.14748e+07 + -3.96754e+06 = 1.75073e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000100110111100000010100011111", b"01001011101000111101001110010010"), -- 2.14748e+07 + -1776.16 = 2.14731e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"01001011101000111101011100001010"), -- 2.14748e+07 + -0.18 = 2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001100001000111101011100001010"), -- -2.14748e+07 + -2.14748e+07 = -4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"01000011001010110000101000111101", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011010110100"), -- 171.04 + -2.14748e+07 = -2.14747e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"01001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001100001000111101011100001010"), -- 2.14748e+07 + 2.14748e+07 = 4.29497e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"11001011101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11001011101000111101011100001010"), -- -2.14748e+07 + 0 = -2.14748e+07
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11001011101000111101011100001010", b"11001011101000111101011100001010"), -- 0 + -2.14748e+07 = -2.14748e+07
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01001011101000111101011100001010", b"01001011101000111101011100001010"), -- -0 + 2.14748e+07 = 2.14748e+07
	(b"11000111110101110111011011000110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000111110101110111011011000110"), -- -110318 + -0 = -110318

	(b"11000001010110100001010001111011", b"00000000000000000000000000000000"),
	(b"11000010001010000001111010111000", b"11000010010111101010001111010111"), -- -13.63 + -42.03 = -55.66
	(b"11000010001111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110001010111010111000011", b"11000011000100011011101011100010"), -- -47 + -98.73 = -145.73
	(b"01000010101000010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001000110011001100110011", b"01000010000111101100110011001101"), -- 80.5 + -40.8 = 39.7
	(b"11000010011111011111010111000011", b"00000000000000000000000000000000"),
	(b"11000010101010101000111101011100", b"11000011000101001100010100011111"), -- -63.49 + -85.28 = -148.77
	(b"01000010000101111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010010100100001111010111000", b"01000010101101001111101011100001"), -- 37.96 + 52.53 = 90.49
	(b"11000010001011101010001111010111", b"00000000000000000000000000000000"),
	(b"01000010010010001110000101001000", b"01000000110100011110101110001000"), -- -43.66 + 50.22 = 6.56
	(b"01000010011010100111000010100100", b"00000000000000000000000000000000"),
	(b"11000001110000000010100011110110", b"01000010000010100101110000101001"), -- 58.61 + -24.02 = 34.59
	(b"11000010010001101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010000011001100110011001101", b"11000001011010001010001111011000"), -- -49.74 + 35.2 = -14.54
	(b"01000001100011111101011100001010", b"00000000000000000000000000000000"),
	(b"11000010100010111111000010100100", b"11000010010011111111010111000011"), -- 17.98 + -69.97 = -51.99
	(b"01000010001111111011100001010010", b"00000000000000000000000000000000"),
	(b"11000010000000001110000101001000", b"01000001011110110101110000101000"), -- 47.93 + -32.22 = 15.71
	(b"11000001101110110111000010100100", b"00000000000000000000000000000000"),
	(b"01000001100010111010111000010100", b"11000000101111110000101001000000"), -- -23.43 + 17.46 = -5.97
	(b"11000010010000100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100000010111000010100100", b"11000010000000010100011110101110"), -- -48.5 + 16.18 = -32.32
	(b"11000010101010010100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100000110000101000111101", b"11000010100010001000101000111110"), -- -84.65 + 16.38 = -68.27
	(b"01000010001110010001010001111011", b"00000000000000000000000000000000"),
	(b"11000010000101111101011100001010", b"01000001000001001111010111000100"), -- 46.27 + -37.96 = 8.31
	(b"01000010101001011101000111101100", b"00000000000000000000000000000000"),
	(b"11000001010101100001010001111011", b"01000010100010110000111101011101"), -- 82.91 + -13.38 = 69.53
	(b"01000010001111011010111000010100", b"00000000000000000000000000000000"),
	(b"11000001110101100111101011100001", b"01000001101001001110000101000111"), -- 47.42 + -26.81 = 20.61
	(b"01000010101000110100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000100001000010100011111", b"01000010001101100001010001111011"), -- 81.65 + -36.13 = 45.52
	(b"11000000111110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000010100001101010111000010100", b"11000010100101100110011001100110"), -- -7.86 + -67.34 = -75.2
	(b"01000010100110110101011100001010", b"00000000000000000000000000000000"),
	(b"11000010000110010001111010111000", b"01000010000111011000111101011100"), -- 77.67 + -38.28 = 39.39
	(b"11000010100111001101110000101001", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"11000010100111011110101110000101"), -- -78.43 + -0.53 = -78.96
	(b"11000010101001111111101011100001", b"00000000000000000000000000000000"),
	(b"11000010010000000100011110101110", b"11000011000001000000111101011100"), -- -83.99 + -48.07 = -132.06
	(b"11000010001110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100101101011100001010010", b"11000001110110101110000101001000"), -- -46.2 + 18.84 = -27.36
	(b"01000010100010010110000101001000", b"00000000000000000000000000000000"),
	(b"01000010000001111111010111000011", b"01000010110011010101110000101010"), -- 68.69 + 33.99 = 102.68
	(b"11000001101100010111000010100100", b"00000000000000000000000000000000"),
	(b"01000010011100010110011001100110", b"01000010000110001010111000010100"), -- -22.18 + 60.35 = 38.17
	(b"01000010100011010001111010111000", b"00000000000000000000000000000000"),
	(b"11000010011111010000101000111101", b"01000000111010011001100110011000"), -- 70.56 + -63.26 = 7.3
	(b"01000001111100010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000110010111101011100001010", b"01000001101111100010100011110110"), -- 30.14 + -6.37 = 23.77
	(b"01000010101100001011100001010010", b"00000000000000000000000000000000"),
	(b"11000010100100011101000111101100", b"01000001011101110011001100110000"), -- 88.36 + -72.91 = 15.45
	(b"11000010101001001010111000010100", b"00000000000000000000000000000000"),
	(b"11000010110001000011001100110011", b"11000011001101000111000010100100"), -- -82.34 + -98.1 = -180.44
	(b"01000010010111011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011010000010100011111", b"01000011000011011111010111000011"), -- 55.45 + 86.51 = 141.96
	(b"01000010011011101111010111000011", b"00000000000000000000000000000000"),
	(b"11000010011010000111000010100100", b"00111111110100001010001111100000"), -- 59.74 + -58.11 = 1.63
	(b"01000010001110111000111101011100", b"00000000000000000000000000000000"),
	(b"01000010101101001000000000000000", b"01000011000010010010001111010111"), -- 46.89 + 90.25 = 137.14
	(b"01000010010101001010111000010100", b"00000000000000000000000000000000"),
	(b"11000001100110000101000111101100", b"01000010000010001000010100011110"), -- 53.17 + -19.04 = 34.13
	(b"01000001101111110111000010100100", b"00000000000000000000000000000000"),
	(b"11000001110101001000111101011100", b"11000000001010001111010111000000"), -- 23.93 + -26.57 = -2.64
	(b"01000010000111100011110101110001", b"00000000000000000000000000000000"),
	(b"01000010001001010011110101110001", b"01000010101000011011110101110001"), -- 39.56 + 41.31 = 80.87
	(b"01000010001111000000101000111101", b"00000000000000000000000000000000"),
	(b"01000001100010001100110011001101", b"01000010100000000011100001010010"), -- 47.01 + 17.1 = 64.11
	(b"10111111101010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000001011111101000111101011100", b"11000001100010011101011100001010"), -- -1.32 + -15.91 = -17.23
	(b"01000010100000100100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000010111101011100001", b"11000001011110010111000010100000"), -- 65.15 + -80.74 = -15.59
	(b"01000010011110101001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101011100001010001111011", b"01000010100000000000010100011111"), -- 62.65 + 1.36 = 64.01
	(b"01000001101001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101010101111010111000011", b"11000010100000010100001010010000"), -- 20.85 + -85.48 = -64.63
	(b"11000010101110011011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100011011101000111101100", b"11000001101011111000010100011100"), -- -92.85 + 70.91 = -21.94
	(b"11000010011100011110000101001000", b"00000000000000000000000000000000"),
	(b"01000001111001110000101000111101", b"11000001111111001011100001010011"), -- -60.47 + 28.88 = -31.59
	(b"11000010000110000011110101110001", b"00000000000000000000000000000000"),
	(b"01000000000101011100001010001111", b"11000010000011101110000101001000"), -- -38.06 + 2.34 = -35.72
	(b"11000010100111010101000111101100", b"00000000000000000000000000000000"),
	(b"01000010110000010000111101011100", b"01000001100011101111010111000000"), -- -78.66 + 96.53 = 17.87
	(b"01000010011001011000010100011111", b"00000000000000000000000000000000"),
	(b"01000001000000110101110000101001", b"01000010100000110010111000010101"), -- 57.38 + 8.21 = 65.59
	(b"01000010001101010111000010100100", b"00000000000000000000000000000000"),
	(b"11000010101101101000111101011100", b"11000010001101111010111000010100"), -- 45.36 + -91.28 = -45.92
	(b"01000010000010001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110000101101011100001010", b"01000011000000111001000111101100"), -- 34.15 + 97.42 = 131.57
	(b"01000010100011000001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001111100011001100110011", b"01000010111010110011001100110100"), -- 70.05 + 47.55 = 117.6
	(b"11000000111100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000010001011111011100001010010", b"11000010010011011100110011001101"), -- -7.52 + -43.93 = -51.45
	(b"01000010101001101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001100011100011110101110001", b"01000010100000110101000111101100"), -- 83.44 + -17.78 = 65.66
	(b"11000010100001110010100011110110", b"00000000000000000000000000000000"),
	(b"11000001111101100111101011100001", b"11000010110001001100011110101110"), -- -67.58 + -30.81 = -98.39
	(b"01000000110011111010111000010100", b"00000000000000000000000000000000"),
	(b"11000001000001110000101000111101", b"10111111111110011001100110011000"), -- 6.49 + -8.44 = -1.95
	(b"01000001101001101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010011101011110000101001000", b"01000010101001001010111000010101"), -- 20.87 + 61.47 = 82.34
	(b"01000001101111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000111100000101000111101100", b"01000001111110100010100011110110"), -- 23.76 + 7.51 = 31.27
	(b"01000010100011100101110000101001", b"00000000000000000000000000000000"),
	(b"11000010010000100001010001111011", b"01000001101101010100011110101110"), -- 71.18 + -48.52 = 22.66
	(b"01000001001101010100011110101110", b"00000000000000000000000000000000"),
	(b"11000001011101001100110011001101", b"11000000011111100001010001111100"), -- 11.33 + -15.3 = -3.97
	(b"01000010100001110101000111101100", b"00000000000000000000000000000000"),
	(b"11000001110000001010001111010111", b"01000010001011100101000111101100"), -- 67.66 + -24.08 = 43.58
	(b"11000010010010011010111000010100", b"00000000000000000000000000000000"),
	(b"01000010010111010011001100110011", b"01000000100111000010100011111000"), -- -50.42 + 55.3 = 4.88
	(b"01000010100100101011110101110001", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"01000010100100101001010001111011"), -- 73.37 + -0.08 = 73.29
	(b"11000001110111000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101001100000101000111101", b"01000010010111011110000101000111"), -- -27.55 + 83.02 = 55.47
	(b"01000010101000111011100001010010", b"00000000000000000000000000000000"),
	(b"11000010100110011010111000010100", b"01000000101000001010001111100000"), -- 81.86 + -76.84 = 5.02
	(b"11000010001011001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000000110111101011100001", b"11000001001001000111101011100100"), -- -43.15 + 32.87 = -10.28
	(b"01000010101001011100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011100001010001111011", b"01000010101010100011110101110001"), -- 82.9 + 2.22 = 85.12
	(b"11000010011110110000101000111101", b"00000000000000000000000000000000"),
	(b"11000001010011110000101000111101", b"11000010100101110110011001100110"), -- -62.76 + -12.94 = -75.7
	(b"01000001111101111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010100111001011100001010010", b"01000010110110101010111000010100"), -- 30.98 + 78.36 = 109.34
	(b"11000010010000001111010111000011", b"00000000000000000000000000000000"),
	(b"11000010011111101110101110000101", b"11000010110111111111000010100100"), -- -48.24 + -63.73 = -111.97
	(b"11000010101110110010100011110110", b"00000000000000000000000000000000"),
	(b"00111111100010100011110101110001", b"11000010101110010000000000000000"), -- -93.58 + 1.08 = -92.5
	(b"11000001100000001011100001010010", b"00000000000000000000000000000000"),
	(b"11000001010011010111000010100100", b"11000001111001110111000010100100"), -- -16.09 + -12.84 = -28.93
	(b"01000010110001110111010111000011", b"00000000000000000000000000000000"),
	(b"01000010101000001011001100110011", b"01000011001101000001010001111011"), -- 99.73 + 80.35 = 180.08
	(b"11000001011110101011100001010010", b"00000000000000000000000000000000"),
	(b"01000001111101000000000000000000", b"01000001011011010100011110101110"), -- -15.67 + 30.5 = 14.83
	(b"11000010011011101001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110011001100110011001101", b"11000010101010101000000000000000"), -- -59.65 + -25.6 = -85.25
	(b"11000010000111110011110101110001", b"00000000000000000000000000000000"),
	(b"11000001000110100011110101110001", b"11000010010001011100110011001101"), -- -39.81 + -9.64 = -49.45
	(b"11000010101000100011100001010010", b"00000000000000000000000000000000"),
	(b"11000001101101001010001111010111", b"11000010110011110110000101001000"), -- -81.11 + -22.58 = -103.69
	(b"11000010000110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011101011110101110000101", b"11000010010101111110000101000111"), -- -38.6 + -15.37 = -53.97
	(b"11000010010001101111010111000011", b"00000000000000000000000000000000"),
	(b"11000001001111010100011110101110", b"11000010011101100100011110101110"), -- -49.74 + -11.83 = -61.57
	(b"10111111101110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000010100011001110000101001000", b"01000010100010011111010111000011"), -- -1.46 + 70.44 = 68.98
	(b"11000010101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001111110100011110101110", b"11000010001110100101000111101100"), -- -94.4 + 47.82 = -46.58
	(b"11000010000001101100001010001111", b"00000000000000000000000000000000"),
	(b"11000010010001010110011001100110", b"11000010101001100001010001111010"), -- -33.69 + -49.35 = -83.04
	(b"01000001011100111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010000101111110101110000101", b"01000010010101001100110011001101"), -- 15.22 + 37.98 = 53.2
	(b"01000010100011000101011100001010", b"00000000000000000000000000000000"),
	(b"11000010101011001100011110101110", b"11000001100000011100001010010000"), -- 70.17 + -86.39 = -16.22
	(b"01000010101101111000111101011100", b"00000000000000000000000000000000"),
	(b"11000001100101011101011100001010", b"01000010100100100001100110011010"), -- 91.78 + -18.73 = 73.05
	(b"11000010101011000100011110101110", b"00000000000000000000000000000000"),
	(b"01000010100001101011110101110001", b"11000001100101100010100011110100"), -- -86.14 + 67.37 = -18.77
	(b"11000010010111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001101011000111101011100", b"11000010110010010010111000010100"), -- -55.2 + -45.39 = -100.59
	(b"11000010101111001010100011110110", b"00000000000000000000000000000000"),
	(b"11000010001110110101000111101100", b"11000011000011010010100011110110"), -- -94.33 + -46.83 = -141.16
	(b"11000001010000111000010100011111", b"00000000000000000000000000000000"),
	(b"01000001101000000001010001111011", b"01000000111110010100011110101110"), -- -12.22 + 20.01 = 7.79
	(b"11000010100000001010100011110110", b"00000000000000000000000000000000"),
	(b"11000000001111110101110000101001", b"11000010100001101010001111010111"), -- -64.33 + -2.99 = -67.32
	(b"01000010011101100111000010100100", b"00000000000000000000000000000000"),
	(b"01000010101011011110101110000101", b"01000011000101001001000111101100"), -- 61.61 + 86.96 = 148.57
	(b"11000010100100011111101011100001", b"00000000000000000000000000000000"),
	(b"01000001111100001000111101011100", b"11000010001010111010111000010100"), -- -72.99 + 30.07 = -42.92
	(b"11000010110001100100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101000011010111000010100", b"11000001100100100111101011100100"), -- -99.15 + 80.84 = -18.31
	(b"11000010100101111100001010001111", b"00000000000000000000000000000000"),
	(b"01000010101010100111000010100100", b"01000001000101010111000010101000"), -- -75.88 + 85.22 = 9.34
	(b"01000010101111100111000010100100", b"00000000000000000000000000000000"),
	(b"01000010101100010010001111010111", b"01000011001101111100101000111110"), -- 95.22 + 88.57 = 183.79
	(b"01000010101111111101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000000001010001111010111", b"01000010110000111101011100001011"), -- 95.91 + 2.01 = 97.92
	(b"11000010100100011000111101011100", b"00000000000000000000000000000000"),
	(b"11000010101001111111000010100100", b"11000011000111001100000000000000"), -- -72.78 + -83.97 = -156.75
	(b"01000010100101110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101011001100011110101110", b"01000011001000011110001111010111"), -- 75.5 + 86.39 = 161.89
	(b"01000001100000000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000100101101011100001010010", b"01000001001101010100011110101111"), -- 16.04 + -4.71 = 11.33
	(b"01000010101100110100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100001111011100001010010", b"01000011000111010111110101110000"), -- 89.63 + 67.86 = 157.49
	(b"01000001101110111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010000000001110101110000101", b"01000010010111101010111000010100"), -- 23.44 + 32.23 = 55.67
	(b"01000010110000100101011100001010", b"00000000000000000000000000000000"),
	(b"11000010100001010110011001100110", b"01000001111100111100001010010000"), -- 97.17 + -66.7 = 30.47
	(b"01000010100000101010111000010100", b"00000000000000000000000000000000"),
	(b"01000010011010101100001010001111", b"01000010111110000000111101011100"), -- 65.34 + 58.69 = 124.03
	(b"01000010101001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101001000110101110000101", b"10111100001000111110000000000000"), -- 82.2 + -82.21 = -0.0100021
	(b"11000010011000110111101011100001", b"00000000000000000000000000000000"),
	(b"11000010100110100001100110011010", b"11000011000001011110101110000101"), -- -56.87 + -77.05 = -133.92
	(b"01000010100111001001100110011010", b"00000000000000000000000000000000"),
	(b"01000001010100101000111101011100", b"01000010101101101110101110000110"), -- 78.3 + 13.16 = 91.46
	(b"11000001101000010000101000111101", b"00000000000000000000000000000000"),
	(b"11000010011011000001111010111000", b"11000010100111100101000111101011"), -- -20.13 + -59.03 = -79.16
	(b"01000010100000011100011110101110", b"00000000000000000000000000000000"),
	(b"01000010010010111111010111000011", b"01000010111001111100001010010000"), -- 64.89 + 50.99 = 115.88
	(b"11000001110101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101111100110011001100110", b"11000010111100110110011001100110"), -- -26.5 + -95.2 = -121.7
	(b"11000001101100100011110101110001", b"00000000000000000000000000000000"),
	(b"01000010101110111111010111000011", b"01000010100011110110011001100111"), -- -22.28 + 93.98 = 71.7
	(b"11000010100001100110000101001000", b"00000000000000000000000000000000"),
	(b"10111111110010111000010100011111", b"11000010100010011000111101011100"), -- -67.19 + -1.59 = -68.78
	(b"01000010101101101010001111010111", b"00000000000000000000000000000000"),
	(b"11000001110111000111101011100001", b"01000010011111110000101000111110"), -- 91.32 + -27.56 = 63.76
	(b"11000001010000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000010100001001000111101011100", b"11000010100111001011100001010010"), -- -12.08 + -66.28 = -78.36
	(b"01000010100101101010001111010111", b"00000000000000000000000000000000"),
	(b"11000010001110011000111101011100", b"01000001111001110111000010100100"), -- 75.32 + -46.39 = 28.93
	(b"11000010100100110100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100100110011110101110001", b"10111100001000111100000000000000"), -- -73.63 + 73.62 = -0.00999451
	(b"00111111100101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000010110001000111101011100001", b"01000010110001101100110011001101"), -- 1.16 + 98.24 = 99.4
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001001010100011110110", b"11000010110001011111010111000011"), -- -0.65 + -98.33 = -98.98
	(b"11000010011110110011110101110001", b"00000000000000000000000000000000"),
	(b"11000010110000111001010001111011", b"11000011001000001001100110011010"), -- -62.81 + -97.79 = -160.6
	(b"01000001110010110111000010100100", b"00000000000000000000000000000000"),
	(b"11000010100101010001100110011010", b"11000010010001000111101011100010"), -- 25.43 + -74.55 = -49.12
	(b"11000000110011111010111000010100", b"00000000000000000000000000000000"),
	(b"11000010101011111110101110000101", b"11000010101111001110011001100110"), -- -6.49 + -87.96 = -94.45
	(b"11000010110000101000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100100111101000111101100", b"11000001101110101011100001010000"), -- -97.25 + 73.91 = -23.34
	(b"01000010010011100101110000101001", b"00000000000000000000000000000000"),
	(b"01000010011111011110000101001000", b"01000010111001100001111010111000"), -- 51.59 + 63.47 = 115.06
	(b"01000001101010110100011110101110", b"00000000000000000000000000000000"),
	(b"01000010000000000011110101110001", b"01000010010101011110000101001000"), -- 21.41 + 32.06 = 53.47
	(b"01000010001100001001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111101001010001111010111", b"01000001010110010001111010111010"), -- 44.15 + -30.58 = 13.57
	(b"01000010011001010101000111101100", b"00000000000000000000000000000000"),
	(b"11000010000011110111000010100100", b"01000001101010111100001010010000"), -- 57.33 + -35.86 = 21.47
	(b"11000010000000000001010001111011", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"11000001111110011101011100001010"), -- -32.02 + 0.79 = -31.23
	(b"11000010011001001010001111010111", b"00000000000000000000000000000000"),
	(b"01000001111011011000010100011111", b"11000001110110111100001010001111"), -- -57.16 + 29.69 = -27.47
	(b"01000010100001011101110000101001", b"00000000000000000000000000000000"),
	(b"01000010010011001010111000010100", b"01000010111011000011001100110011"), -- 66.93 + 51.17 = 118.1
	(b"11000001011001110000101000111101", b"00000000000000000000000000000000"),
	(b"01000010100000100111010111000011", b"01000010010010110010100011110111"), -- -14.44 + 65.23 = 50.79
	(b"11000001110110111110101110000101", b"00000000000000000000000000000000"),
	(b"01000010000111010111101011100001", b"01000001001111100001010001111010"), -- -27.49 + 39.37 = 11.88
	(b"01000010001100110100011110101110", b"00000000000000000000000000000000"),
	(b"01000010100110000111000010100100", b"01000010111100100001010001111011"), -- 44.82 + 76.22 = 121.04
	(b"11000010110000111101110000101001", b"00000000000000000000000000000000"),
	(b"11000010100000101010100011110110", b"11000011001000110100001010010000"), -- -97.93 + -65.33 = -163.26
	(b"01000010101000011111000010100100", b"00000000000000000000000000000000"),
	(b"11000010101101111111010111000011", b"11000001001100000010100011111000"), -- 80.97 + -91.98 = -11.01
	(b"01000010010111001111010111000011", b"00000000000000000000000000000000"),
	(b"11000001111101101010001111010111", b"01000001110000110100011110101111"), -- 55.24 + -30.83 = 24.41
	(b"01000010100111101111010111000011", b"00000000000000000000000000000000"),
	(b"11000010010111000111101011100001", b"01000001110000101110000101001010"), -- 79.48 + -55.12 = 24.36
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001011100111101011100001", b"01000010000111110100011110101110"), -- -3.8 + 43.62 = 39.82
	(b"01000001011011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110101110000101000111101", b"01000010001001110001111010111000"), -- 14.9 + 26.88 = 41.78
	(b"11000010010100110000101000111101", b"00000000000000000000000000000000"),
	(b"11000010011011001010111000010100", b"11000010110111111101110000101000"), -- -52.76 + -59.17 = -111.93
	(b"11000010100101010111101011100001", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"11000010100101101011001100110011"), -- -74.74 + -0.61 = -75.35
	(b"01000010000101001110101110000101", b"00000000000000000000000000000000"),
	(b"01000010000010010101110000101001", b"01000010100011110010001111010111"), -- 37.23 + 34.34 = 71.57
	(b"01000000111110101000111101011100", b"00000000000000000000000000000000"),
	(b"01000010001111110011001100110011", b"01000010010111101000010100011110"), -- 7.83 + 47.8 = 55.63
	(b"01000001100000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001111111000110011001100110", b"01000010001111100110011001100110"), -- 16.05 + 31.55 = 47.6
	(b"00111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000010010100100010100011110110", b"11000010010100100000101000111110"), -- 0.03 + -52.54 = -52.51
	(b"11000000111010001010001111010111", b"00000000000000000000000000000000"),
	(b"11000010011010111000111101011100", b"11000010100001000101000111101011"), -- -7.27 + -58.89 = -66.16
	(b"11000001001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110001100100011110101110", b"11000010110110100100011110101110"), -- -10 + -99.14 = -109.14
	(b"11000001100111010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101100101010111000010100", b"11000010110110011111101011100001"), -- -19.65 + -89.34 = -108.99
	(b"01000010100101010100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011001010111101011100001", b"01000001100010100011110101110010"), -- 74.65 + -57.37 = 17.28
	(b"11000010000111010000101000111101", b"00000000000000000000000000000000"),
	(b"11000001010101001010001111010111", b"11000010010100100011001100110011"), -- -39.26 + -13.29 = -52.55
	(b"11000010010101001000010100011111", b"00000000000000000000000000000000"),
	(b"11000010101101101011100001010010", b"11000011000100000111110101110001"), -- -53.13 + -91.36 = -144.49
	(b"11000010101010001101110000101001", b"00000000000000000000000000000000"),
	(b"11000010100101000111010111000011", b"11000011000111101010100011110110"), -- -84.43 + -74.23 = -158.66
	(b"01000001100011010111000010100100", b"00000000000000000000000000000000"),
	(b"01000010001100110110011001100110", b"01000010011110100001111010111000"), -- 17.68 + 44.85 = 62.53
	(b"11000010010110101000010100011111", b"00000000000000000000000000000000"),
	(b"01000000110000000101000111101100", b"11000010010000100111101011100010"), -- -54.63 + 6.01 = -48.62
	(b"11000001110110100000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101001100001010001111011", b"11000010000000011100001010001111"), -- -27.25 + -5.19 = -32.44
	(b"11000010101101011111010111000011", b"00000000000000000000000000000000"),
	(b"01000001010100111101011100001010", b"11000010100110110111101011100010"), -- -90.98 + 13.24 = -77.74
	(b"11000000110010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000010110000101101011100001010", b"01000010101101100010100011110110"), -- -6.34 + 97.42 = 91.08
	(b"01000001010101011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010100000101001100110011010", b"01000010100111010101011100001011"), -- 13.37 + 65.3 = 78.67
	(b"01000010001000000101110000101001", b"00000000000000000000000000000000"),
	(b"11000010100101110110101110000101", b"11000010000011100111101011100001"), -- 40.09 + -75.71 = -35.62
	(b"11000010101100110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110111100111101011100001", b"11000010111010110000010100011110"), -- -89.7 + -27.81 = -117.51
	(b"01000001100010100001010001111011", b"00000000000000000000000000000000"),
	(b"01000010100011111101000111101100", b"01000010101100100101011100001011"), -- 17.26 + 71.91 = 89.17
	(b"01000010110000000100001010001111", b"00000000000000000000000000000000"),
	(b"01000010110001110001111010111000", b"01000011010000111011000010100100"), -- 96.13 + 99.56 = 195.69
	(b"01000010101011110001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101001000010111000010100", b"01000000101011101011100001100000"), -- 87.55 + -82.09 = 5.46001
	(b"01000010010011111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010001101011101011100001010", b"01000010110000101010111000010100"), -- 51.88 + 45.46 = 97.34
	(b"01000010100000001000101000111101", b"00000000000000000000000000000000"),
	(b"11000010010010111111010111000011", b"01000001010101000111101011011100"), -- 64.27 + -50.99 = 13.28
	(b"11000010010100101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010010111110101000111101100", b"01000000010001011100001010010000"), -- -52.74 + 55.83 = 3.09
	(b"11000001111001100011110101110001", b"00000000000000000000000000000000"),
	(b"11000010100101000010100011110110", b"11000010110011011011100001010010"), -- -28.78 + -74.08 = -102.86
	(b"01000001110001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010110110011001100110011", b"11000001111100000110011001100110"), -- 24.75 + -54.8 = -30.05
	(b"11000010100101111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101100110001100110011010", b"01000001010111000000000000000000"), -- -75.8 + 89.55 = 13.75
	(b"11000010011110000001010001111011", b"00000000000000000000000000000000"),
	(b"00111111110011110101110000101001", b"11000010011100011001100110011010"), -- -62.02 + 1.62 = -60.4
	(b"01000010101001011001111010111000", b"00000000000000000000000000000000"),
	(b"11000010010010011000111101011100", b"01000010000000011010111000010100"), -- 82.81 + -50.39 = 32.42
	(b"11000010000001101000010100011111", b"00000000000000000000000000000000"),
	(b"11000010010011011000111101011100", b"11000010101010100000101000111110"), -- -33.63 + -51.39 = -85.02
	(b"11000001111000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101101110111010111000011", b"01000010011111100001111010111001"), -- -28.2 + 91.73 = 63.53
	(b"11000010000011110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100010110101000111101100", b"11000010110100101101000111101100"), -- -35.75 + -69.66 = -105.41
	(b"01000001100011110001111010111000", b"00000000000000000000000000000000"),
	(b"01000001100001001111010111000011", b"01000010000010100000101000111110"), -- 17.89 + 16.62 = 34.51
	(b"11000010101111001011110101110001", b"00000000000000000000000000000000"),
	(b"01000010100111010100011110101110", b"11000001011110111010111000011000"), -- -94.37 + 78.64 = -15.73
	(b"01000010011111001011100001010010", b"00000000000000000000000000000000"),
	(b"01000001011001110011001100110011", b"01000010100110110100001010001111"), -- 63.18 + 14.45 = 77.63
	(b"11000001101000101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001100100101111010111000011", b"11000010000110101110101110000110"), -- -20.36 + -18.37 = -38.73
	(b"01000010101111001101000111101100", b"00000000000000000000000000000000"),
	(b"11000010011110010010100011110110", b"01000010000000000111101011100010"), -- 94.41 + -62.29 = 32.12
	(b"11000010100110010001111010111000", b"00000000000000000000000000000000"),
	(b"11000010100000011000000000000000", b"11000011000011010100111101011100"), -- -76.56 + -64.75 = -141.31
	(b"01000010101010010110101110000101", b"00000000000000000000000000000000"),
	(b"01000001001101000101000111101100", b"01000010101111111111010111000010"), -- 84.71 + 11.27 = 95.98
	(b"11000010101000101000101000111101", b"00000000000000000000000000000000"),
	(b"11000010010101001101011100001010", b"11000011000001100111101011100001"), -- -81.27 + -53.21 = -134.48
	(b"01000010000011100000101000111101", b"00000000000000000000000000000000"),
	(b"01000010101101011111101011100001", b"01000010111111010000000000000000"), -- 35.51 + 90.99 = 126.5
	(b"11000010011000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100000101111010111000011", b"01000001000010010100011110110000"), -- -56.9 + 65.48 = 8.58
	(b"11000010010001110010100011110110", b"00000000000000000000000000000000"),
	(b"01000010110001001100110011001101", b"01000010010000100111000010100100"), -- -49.79 + 98.4 = 48.61
	(b"01000010001110000011110101110001", b"00000000000000000000000000000000"),
	(b"01000010000000101000010100011111", b"01000010100111010110000101001000"), -- 46.06 + 32.63 = 78.69
	(b"01000001111111001010001111010111", b"00000000000000000000000000000000"),
	(b"11000010100010001111101011100001", b"11000010000100111010001111010110"), -- 31.58 + -68.49 = -36.91
	(b"01000001110111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001111000000000000000", b"01000010110111110110011001100110"), -- 27.95 + 83.75 = 111.7
	(b"11000001110011000111101011100001", b"00000000000000000000000000000000"),
	(b"01000010100101100110000101001000", b"01000010010001101000010100100000"), -- -25.56 + 75.19 = 49.63
	(b"01000010001101011010001111010111", b"00000000000000000000000000000000"),
	(b"11000010101111101111101011100001", b"11000010010010000101000111101011"), -- 45.41 + -95.49 = -50.08
	(b"11000001000001010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010101011110011001100110011", b"01000010100111101000101000111101"), -- -8.33 + 87.6 = 79.27
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010011011010001111010111", b"01000010010101110011110101110001"), -- 2.4 + 51.41 = 53.81
	(b"11000010001000011000010100011111", b"00000000000000000000000000000000"),
	(b"01000001101011011001100110011010", b"11000001100101010111000010100100"), -- -40.38 + 21.7 = -18.68
	(b"01000001111110101000111101011100", b"00000000000000000000000000000000"),
	(b"01000010100100000100110011001101", b"01000010110011101111000010100100"), -- 31.32 + 72.15 = 103.47
	(b"01000010101001000011100001010010", b"00000000000000000000000000000000"),
	(b"11000010000010011011100001010010", b"01000010001111101011100001010010"), -- 82.11 + -34.43 = 47.68
	(b"11000001100110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100100100101110000101001", b"11000010101110000111010111000010"), -- -19.05 + -73.18 = -92.23
	(b"01000010100110011100001010001111", b"00000000000000000000000000000000"),
	(b"11000001011001111000010100011111", b"01000010011110011010001111010110"), -- 76.88 + -14.47 = 62.41
	(b"01000010010111001101011100001010", b"00000000000000000000000000000000"),
	(b"01000010000001111011100001010010", b"01000010101100100100011110101110"), -- 55.21 + 33.93 = 89.14
	(b"11000001100111010101110000101001", b"00000000000000000000000000000000"),
	(b"01000010100111000110000101001000", b"01000010011010100001010001111100"), -- -19.67 + 78.19 = 58.52
	(b"01000010001110000011110101110001", b"00000000000000000000000000000000"),
	(b"01000010001000100111000010100100", b"01000010101011010101011100001010"), -- 46.06 + 40.61 = 86.67
	(b"11000010100100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000110111111010111000011", b"11000010000010110011110101110001"), -- -73.8 + 38.99 = -34.81
	(b"01000010000100011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101100000111101011100001", b"11000010010011110010100011110101"), -- 36.45 + -88.24 = -51.79
	(b"11000001101111000011110101110001", b"00000000000000000000000000000000"),
	(b"01000000011100011110101110000101", b"11000001100111100000000000000000"), -- -23.53 + 3.78 = -19.75
	(b"01000010101111000100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101100011100001010001111", b"01000000101010001010001111100000"), -- 94.15 + -88.88 = 5.27
	(b"01000010101111100001111010111000", b"00000000000000000000000000000000"),
	(b"01000010000010111010001111010111", b"01000011000000011111100001010010"), -- 95.06 + 34.91 = 129.97
	(b"01000010011110011100001010001111", b"00000000000000000000000000000000"),
	(b"11000010100011111110011001100110", b"11000001000110000010100011110100"), -- 62.44 + -71.95 = -9.51
	(b"11000010000111010101110000101001", b"00000000000000000000000000000000"),
	(b"10111111100001010001111010111000", b"11000010001000011000010100011111"), -- -39.34 + -1.04 = -40.38
	(b"10111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000010100000000101000111101100", b"11000010100000001000111101011101"), -- -0.12 + -64.16 = -64.28
	(b"11000010100100100101011100001010", b"00000000000000000000000000000000"),
	(b"11000010001000111000111101011100", b"11000010111001000001111010111000"), -- -73.17 + -40.89 = -114.06
	(b"01000001100011011100001010001111", b"00000000000000000000000000000000"),
	(b"11000001111110101111010111000011", b"11000001010110100110011001101000"), -- 17.72 + -31.37 = -13.65
	(b"01000010100001000101110000101001", b"00000000000000000000000000000000"),
	(b"01000010001000011100110011001101", b"01000010110101010100001010010000"), -- 66.18 + 40.45 = 106.63
	(b"11000010101111000011100001010010", b"00000000000000000000000000000000"),
	(b"01000010100010000100011110101110", b"11000001110011111100001010010000"), -- -94.11 + 68.14 = -25.97
	(b"11000010011101001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010101100111010111000010100", b"01000001111001011001100110011000"), -- -61.14 + 89.84 = 28.7
	(b"11000010100111111111101011100001", b"00000000000000000000000000000000"),
	(b"11000010100001100011001100110011", b"11000011000100110001011100001010"), -- -79.99 + -67.1 = -147.09
	(b"11000010100000111011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100100011110000101001000", b"01000000111000101110000101010000"), -- -65.85 + 72.94 = 7.09
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001100000010101110000101001", b"11000001100001010100011110101110"), -- -0.49 + -16.17 = -16.66
	(b"01000001111100100001010001111011", b"00000000000000000000000000000000"),
	(b"01000010110001110000000000000000", b"01000011000000011100001010001111"), -- 30.26 + 99.5 = 129.76
	(b"01000001111110100011110101110001", b"00000000000000000000000000000000"),
	(b"01000010011100100011001100110011", b"01000010101101111010100011110110"), -- 31.28 + 60.55 = 91.83
	(b"11000001001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011010001010001111010111", b"01000010001111000011110101110000"), -- -11.1 + 58.16 = 47.06
	(b"01000001101101110001111010111000", b"00000000000000000000000000000000"),
	(b"01000010010011101110101110000101", b"01000010100101010011110101110000"), -- 22.89 + 51.73 = 74.62
	(b"01000000110111011100001010001111", b"00000000000000000000000000000000"),
	(b"11000010101101001001111010111000", b"11000010101001101100001010001111"), -- 6.93 + -90.31 = -83.38
	(b"11000001100011111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010101000010100011111", b"01000010100001101001111010111000"), -- -17.95 + 85.26 = 67.31
	(b"11000010011000110011110101110001", b"00000000000000000000000000000000"),
	(b"11000010100111100101000111101100", b"11000011000001111111100001010010"), -- -56.81 + -79.16 = -135.97
	(b"11000010000110111100001010001111", b"00000000000000000000000000000000"),
	(b"11000000001111100001010001111011", b"11000010001001111010001111010111"), -- -38.94 + -2.97 = -41.91
	(b"01000000101111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000001010000100001010001111011", b"01000001100100001000111101011100"), -- 5.94 + 12.13 = 18.07
	(b"11000010100010101010100011110110", b"00000000000000000000000000000000"),
	(b"11000010100100100100001010001111", b"11000011000011100111010111000010"), -- -69.33 + -73.13 = -142.46
	(b"11000010100001000110101110000101", b"00000000000000000000000000000000"),
	(b"10111111111100011110101110000101", b"11000010100010000011001100110011"), -- -66.21 + -1.89 = -68.1
	(b"11000010001010001110101110000101", b"00000000000000000000000000000000"),
	(b"11000001001011110011001100110011", b"11000010010101001011100001010010"), -- -42.23 + -10.95 = -53.18
	(b"01000010011011011100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110100010011001100110011", b"01000010101010110011001100110011"), -- 59.45 + 26.15 = 85.6
	(b"01000010100111010001111010111000", b"00000000000000000000000000000000"),
	(b"11000001110110000101000111101100", b"01000010010011100001010001111010"), -- 78.56 + -27.04 = 51.52
	(b"01000001100110111100001010001111", b"00000000000000000000000000000000"),
	(b"11000010101111110111101011100001", b"11000010100110001000101000111101"), -- 19.47 + -95.74 = -76.27
	(b"11000010011010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000010101100110011001100110", b"11000010011110001110101110000101"), -- -58.88 + -3.35 = -62.23
	(b"11000001000101111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010011000111100001010001111", b"01000010001111011110000101000111"), -- -9.47 + 56.94 = 47.47
	(b"01000010100010000101110000101001", b"00000000000000000000000000000000"),
	(b"11000001000100010001111010111000", b"01000010011011000111000010100100"), -- 68.18 + -9.07 = 59.11
	(b"01000010101011110111101011100001", b"00000000000000000000000000000000"),
	(b"11000001110101111001100110011010", b"01000010011100110010100011110101"), -- 87.74 + -26.95 = 60.79
	(b"11000010001011111000111101011100", b"00000000000000000000000000000000"),
	(b"11000001000011111101011100001010", b"11000010010100111000010100011110"), -- -43.89 + -8.99 = -52.88
	(b"11000001111010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000010101100100011110101110001", b"11000010111011010001111010111001"), -- -29.44 + -89.12 = -118.56
	(b"11000001111110101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010010011011111010111000011", b"01000001101000001111010111000011"), -- -31.37 + 51.49 = 20.12
	(b"11000010101011001011110101110001", b"00000000000000000000000000000000"),
	(b"11000001011100101000111101011100", b"11000010110010110000111101011100"), -- -86.37 + -15.16 = -101.53
	(b"01000000110101101011100001010010", b"00000000000000000000000000000000"),
	(b"01000010101001110111101011100001", b"01000010101101001110011001100110"), -- 6.71 + 83.74 = 90.45
	(b"11000010101010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101101001101011100001010", b"01000000110011010111000010100000"), -- -84 + 90.42 = 6.42
	(b"01000001100001110111000010100100", b"00000000000000000000000000000000"),
	(b"01000010001101101011100001010010", b"01000010011110100111000010100100"), -- 16.93 + 45.68 = 62.61
	(b"01000001101111000101000111101100", b"00000000000000000000000000000000"),
	(b"11000010101001001110000101001000", b"11000010011010111001100110011010"), -- 23.54 + -82.44 = -58.9
	(b"01000010101000010011110101110001", b"00000000000000000000000000000000"),
	(b"10111111111111010111000010100100", b"01000010100111010100011110101110"), -- 80.62 + -1.98 = 78.64
	(b"11000010101101100001111010111000", b"00000000000000000000000000000000"),
	(b"11000010110000001110101110000101", b"11000011001110111000010100011110"), -- -91.06 + -96.46 = -187.52
	(b"11000010100011000010001111010111", b"00000000000000000000000000000000"),
	(b"11000001101000111010111000010100", b"11000010101101010000111101011100"), -- -70.07 + -20.46 = -90.53
	(b"11000010100101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100110110010100011110110", b"11000011000110001001010001111011"), -- -75 + -77.58 = -152.58
	(b"01000010100111111011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110001101011100001010010", b"01000010010111000000101000111101"), -- 79.85 + -24.84 = 55.01
	(b"01000010100111000000101000111101", b"00000000000000000000000000000000"),
	(b"00111111111001010001111010111000", b"01000010100111111001111010111000"), -- 78.02 + 1.79 = 79.81
	(b"01000010011011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000000010101000111101100", b"01000010101110000100001010010000"), -- 59.8 + 32.33 = 92.13
	(b"01000010100111110100011110101110", b"00000000000000000000000000000000"),
	(b"11000010101000000110000101001000", b"10111111000011001100110100000000"), -- 79.64 + -80.19 = -0.550003
	(b"11000010011110110011110101110001", b"00000000000000000000000000000000"),
	(b"01000010100000011010100011110110", b"01000000000000010100011110110000"), -- -62.81 + 64.83 = 2.02
	(b"01000001111100100101000111101100", b"00000000000000000000000000000000"),
	(b"01000001000110000010100011110110", b"01000010000111110011001100110100"), -- 30.29 + 9.51 = 39.8
	(b"01000001100001011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010101111110110011001100110", b"11000010100111011110101110000101"), -- 16.74 + -95.7 = -78.96
	(b"11000010100010001000010100011111", b"00000000000000000000000000000000"),
	(b"11000010101101101101011100001010", b"11000011000111111010111000010100"), -- -68.26 + -91.42 = -159.68
	(b"11000001010000111000010100011111", b"00000000000000000000000000000000"),
	(b"11000001011000100011110101110001", b"11000001110100101110000101001000"), -- -12.22 + -14.14 = -26.36
	(b"01000010101010110101000111101100", b"00000000000000000000000000000000"),
	(b"11000010000100001000111101011100", b"01000010010001100001010001111100"), -- 85.66 + -36.14 = 49.52
	(b"11000000111010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001101011010001111010111", b"11000010010100101010001111010111"), -- -7.25 + -45.41 = -52.66
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000010101010111110000101001000", b"01000010101011001110101110000101"), -- 0.52 + 85.94 = 86.46
	(b"01000001110111000111101011100001", b"00000000000000000000000000000000"),
	(b"01000010101101011100110011001101", b"01000010111011001110101110000101"), -- 27.56 + 90.9 = 118.46
	(b"11000010110000110010111000010100", b"00000000000000000000000000000000"),
	(b"11000000100000010100011110101110", b"11000010110010110100001010001111"), -- -97.59 + -4.04 = -101.63
	(b"11000010000001110101000111101100", b"00000000000000000000000000000000"),
	(b"01000000111001001100110011001101", b"11000001110101010111000010100101"), -- -33.83 + 7.15 = -26.68
	(b"01000010100011001000101000111101", b"00000000000000000000000000000000"),
	(b"11000010011010101000111101011100", b"01000001001110100001010001111000"), -- 70.27 + -58.64 = 11.63
	(b"01000010101111011000111101011100", b"00000000000000000000000000000000"),
	(b"01000010000000110000101000111101", b"01000010111111110001010001111010"), -- 94.78 + 32.76 = 127.54
	(b"11000010100010101011110101110001", b"00000000000000000000000000000000"),
	(b"01000010001011111110101110000101", b"11000001110010110001111010111010"), -- -69.37 + 43.98 = -25.39
	(b"11000000110100101000111101011100", b"00000000000000000000000000000000"),
	(b"11000010101110001011100001010010", b"11000010110001011110000101001000"), -- -6.58 + -92.36 = -98.94
	(b"01000001101000010111000010100100", b"00000000000000000000000000000000"),
	(b"01000010100100100101110000101001", b"01000010101110101011100001010010"), -- 20.18 + 73.18 = 93.36
	(b"01000010011111000111000010100100", b"00000000000000000000000000000000"),
	(b"01000001100011111010111000010100", b"01000010101000100010001111010111"), -- 63.11 + 17.96 = 81.07
	(b"11000001111110100111101011100001", b"00000000000000000000000000000000"),
	(b"01000010101110001101110000101001", b"01000010011101000111101011100010"), -- -31.31 + 92.43 = 61.12
	(b"01000010000111010011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101001000111101011100001", b"01000010000010001010001111010111"), -- 39.3 + -5.14 = 34.16
	(b"11000001101111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000010100011011000101000111101", b"11000010101111010000111101011100"), -- -23.76 + -70.77 = -94.53
	(b"11000010101010100001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010000010010100011110110", b"11000010000100110000101000111110"), -- -85.05 + 48.29 = -36.76
	(b"01000010100000100001111010111000", b"00000000000000000000000000000000"),
	(b"01000000100100011001100110011010", b"01000010100010110011100001010010"), -- 65.06 + 4.55 = 69.61
	(b"11000010101001001011110101110001", b"00000000000000000000000000000000"),
	(b"11000001101000100001010001111011", b"11000010110011010100001010010000"), -- -82.37 + -20.26 = -102.63
	(b"01000010100100100101011100001010", b"00000000000000000000000000000000"),
	(b"11000010101000000011001100110011", b"11000000110111011100001010010000"), -- 73.17 + -80.1 = -6.93
	(b"01000001101100111110101110000101", b"00000000000000000000000000000000"),
	(b"11000001010101101000111101011100", b"01000001000100010100011110101110"), -- 22.49 + -13.41 = 9.08
	(b"11000010010100010101000111101100", b"00000000000000000000000000000000"),
	(b"01000010011101101000010100011111", b"01000001000101001100110011001100"), -- -52.33 + 61.63 = 9.3
	(b"11000010101101000101011100001010", b"00000000000000000000000000000000"),
	(b"11000001010010010111000010100100", b"11000010110011011000010100011110"), -- -90.17 + -12.59 = -102.76
	(b"11000001001100010111000010100100", b"00000000000000000000000000000000"),
	(b"01000001100101001010001111010111", b"01000000111011111010111000010100"), -- -11.09 + 18.58 = 7.49
	(b"01000010001011111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101110010000000000000000", b"01000011000010000110011001100110"), -- 43.9 + 92.5 = 136.4
	(b"11000010100011110010100011110110", b"00000000000000000000000000000000"),
	(b"01000001100100000010100011110110", b"11000010010101100011110101110001"), -- -71.58 + 18.02 = -53.56
	(b"11000010011011001000010100011111", b"00000000000000000000000000000000"),
	(b"01000010100001100000111101011100", b"01000000111111001100110011001000"), -- -59.13 + 67.03 = 7.9
	(b"11000010001000101000010100011111", b"00000000000000000000000000000000"),
	(b"01000001010110110101110000101001", b"11000001110101110101110000101010"), -- -40.63 + 13.71 = -26.92
	(b"01000010101001110001111010111000", b"00000000000000000000000000000000"),
	(b"11000010101100011010100011110110", b"11000000101010001010001111100000"), -- 83.56 + -88.83 = -5.27
	(b"01000010001111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000100000111101011100001010", b"01000010001010111010111000010101"), -- 47.04 + -4.12 = 42.92
	(b"01000001000001111000010100011111", b"00000000000000000000000000000000"),
	(b"01000001000000101110000101001000", b"01000001100001010011001100110100"), -- 8.47 + 8.18 = 16.65
	(b"01000010101011011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010100111000000000000000000", b"01000001000011110101110000101000"), -- 86.96 + -78 = 8.96
	(b"11000010101100100010100011110110", b"00000000000000000000000000000000"),
	(b"01000010100010111100001010001111", b"11000001100110011001100110011100"), -- -89.08 + 69.88 = -19.2
	(b"11000010100100100111000010100100", b"00000000000000000000000000000000"),
	(b"11000010100100010110000101001000", b"11000011000100011110100011110110"), -- -73.22 + -72.69 = -145.91
	(b"11000000100100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010100100001110011001100110", b"01000010100001111010100011110101"), -- -4.62 + 72.45 = 67.83
	(b"11000001110011010101110000101001", b"00000000000000000000000000000000"),
	(b"01000010010010101010001111010111", b"01000001110001111110101110000101"), -- -25.67 + 50.66 = 24.99
	(b"01000010011001000111000010100100", b"00000000000000000000000000000000"),
	(b"01000010110000110000000000000000", b"01000011000110101001110000101001"), -- 57.11 + 97.5 = 154.61
	(b"11000010000110010000101000111101", b"00000000000000000000000000000000"),
	(b"01000010101001011000010100011111", b"01000010001100100000000000000001"), -- -38.26 + 82.76 = 44.5
	(b"01000010010111001100001010001111", b"00000000000000000000000000000000"),
	(b"01000010010100101000010100011111", b"01000010110101111010001111010111"), -- 55.19 + 52.63 = 107.82
	(b"01000010101101010100001010001111", b"00000000000000000000000000000000"),
	(b"00111111001100001010001111010111", b"01000010101101101010001111010111"), -- 90.63 + 0.69 = 91.32
	(b"01000010100011110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000100100100011110101110", b"01000010000011001000010100011110"), -- 71.7 + -36.57 = 35.13
	(b"11000010101100001010111000010100", b"00000000000000000000000000000000"),
	(b"01000010101111000010001111010111", b"01000000101101110101110000110000"), -- -88.34 + 94.07 = 5.73
	(b"01000001110011001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010110000001001111010111000", b"01000010111100111100001010001111"), -- 25.57 + 96.31 = 121.88
	(b"11000010101110001101000111101100", b"00000000000000000000000000000000"),
	(b"11000010001001100111000010100100", b"11000011000001100000010100011111"), -- -92.41 + -41.61 = -134.02
	(b"11000010100111000101110000101001", b"00000000000000000000000000000000"),
	(b"01000010100100101110011001100110", b"11000000100101110101110000110000"), -- -78.18 + 73.45 = -4.73
	(b"01000010011110110100011110101110", b"00000000000000000000000000000000"),
	(b"11000010000100111010111000010100", b"01000001110011110011001100110100"), -- 62.82 + -36.92 = 25.9
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100111101001100110011010", b"01000010101001010110011001100111"), -- 3.4 + 79.3 = 82.7
	(b"11000010001110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000001101011001000111101011100", b"11000001110010010011001100110100"), -- -46.72 + 21.57 = -25.15
	(b"01000010100101001001010001111011", b"00000000000000000000000000000000"),
	(b"01000010100101010111101011100001", b"01000011000101010000011110101110"), -- 74.29 + 74.74 = 149.03
	(b"11000000110101010001111010111000", b"00000000000000000000000000000000"),
	(b"11000001010001010100011110101110", b"11000001100101111110101110000101"), -- -6.66 + -12.33 = -18.99
	(b"11000010110000111111000010100100", b"00000000000000000000000000000000"),
	(b"11000010101101011000111101011100", b"11000011001111001100000000000000"), -- -97.97 + -90.78 = -188.75
	(b"11000010110000000101110000101001", b"00000000000000000000000000000000"),
	(b"01000010001101100000101000111101", b"11000010010010101010111000010101"), -- -96.18 + 45.51 = -50.67
	(b"01000010101110111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000001010000101000111101100", b"01000010101101101001010001111011"), -- 93.92 + -2.63 = 91.29
	(b"11000010100101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100100010010111000010100", b"11000000010000001010001111100000"), -- -75.6 + 72.59 = -3.01
	(b"01000010010110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010110000000011100001010010", b"01000011000101101110100011110110"), -- 54.8 + 96.11 = 150.91
	(b"11000000100001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000010000001100000101000111101", b"11000010000101101110101110000101"), -- -4.22 + -33.51 = -37.73
	(b"11000010101000100110000101001000", b"00000000000000000000000000000000"),
	(b"01000001111100110001111010111000", b"11000010010010110011001100110100"), -- -81.19 + 30.39 = -50.8
	(b"01000010101001110000010100011111", b"00000000000000000000000000000000"),
	(b"01000010100011011010001111010111", b"01000011000110100101010001111011"), -- 83.51 + 70.82 = 154.33
	(b"11000001100000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101100101000000000000000", b"01000010100100100001100110011010"), -- -16.2 + 89.25 = 73.05
	(b"11000010100001001000101000111101", b"00000000000000000000000000000000"),
	(b"11000001100000000110011001100110", b"11000010101001001010001111010110"), -- -66.27 + -16.05 = -82.32
	(b"11000001101011001110000101001000", b"00000000000000000000000000000000"),
	(b"11000010001110110111000010100100", b"11000010100010001111000010100100"), -- -21.61 + -46.86 = -68.47
	(b"01000010001001110111000010100100", b"00000000000000000000000000000000"),
	(b"11000001000111111000010100011111", b"01000001111111110001111010111000"), -- 41.86 + -9.97 = 31.89
	(b"01000010110000100001111010111000", b"00000000000000000000000000000000"),
	(b"11000001010110101110000101001000", b"01000010101001101100001010001111"), -- 97.06 + -13.68 = 83.38
	(b"01000010101100010101110000101001", b"00000000000000000000000000000000"),
	(b"01000001101010011001100110011010", b"01000010110110111100001010010000"), -- 88.68 + 21.2 = 109.88
	(b"01000000010001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000010100100110111000010100100", b"11000010100011010011100001010010"), -- 3.11 + -73.72 = -70.61
	(b"01000010010011110010100011110110", b"00000000000000000000000000000000"),
	(b"01000010000110010111101011100001", b"01000010101101000101000111101100"), -- 51.79 + 38.37 = 90.16
	(b"11000010001000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101101101010001111010111", b"11000001100011110101110000101001"), -- -40.75 + 22.83 = -17.92
	(b"01000001010101000010100011110110", b"00000000000000000000000000000000"),
	(b"01000010101001001010001111010111", b"01000010101111110010100011110110"), -- 13.26 + 82.32 = 95.58
	(b"01000010000100110000101000111101", b"00000000000000000000000000000000"),
	(b"01000010011000010100011110101110", b"01000010101110100010100011110110"), -- 36.76 + 56.32 = 93.08
	(b"01000001110001100011110101110001", b"00000000000000000000000000000000"),
	(b"11000010100001011110101110000101", b"11000010001010001011100001010010"), -- 24.78 + -66.96 = -42.18
	(b"11000010110001011000111101011100", b"00000000000000000000000000000000"),
	(b"11000010000110001001100110011010", b"11000011000010001110111000010100"), -- -98.78 + -38.15 = -136.93
	(b"11000010101000000100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100100010111101011100001", b"11000000111011000111101011100000"), -- -80.13 + 72.74 = -7.39
	(b"01000010110001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010011000100011110101110", b"01000010001111100001111010111000"), -- 98.6 + -51.07 = 47.53
	(b"01000010011111111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100111111100001010001111", b"01000011000011111101010001111011"), -- 63.95 + 79.88 = 143.83
	(b"01000001101111000011110101110001", b"00000000000000000000000000000000"),
	(b"11000001110011001000111101011100", b"11000000000000101000111101011000"), -- 23.53 + -25.57 = -2.04
	(b"01000010010011011110000101001000", b"00000000000000000000000000000000"),
	(b"11000010101001000001010001111011", b"11000001111101001000111101011100"), -- 51.47 + -82.04 = -30.57
	(b"01000001101001111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010101110000010100011110110", b"01000010111000100000101000111110"), -- 20.94 + 92.08 = 113.02
	(b"11000010101101011000111101011100", b"00000000000000000000000000000000"),
	(b"11000010011111001100110011001101", b"11000011000110011111101011100001"), -- -90.78 + -63.2 = -153.98
	(b"11000001101001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011001110101110000101001", b"01000010000101010101110000101001"), -- -20.5 + 57.84 = 37.34
	(b"11000001110010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110000100011110101110", b"01000010010010110101110000101001"), -- -25.3 + 76.14 = 50.84
	(b"11000010101110011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010001110101110000101001000", b"11000010001110001111010111000010"), -- -92.96 + 46.72 = -46.24
	(b"11000010011111001010111000010100", b"00000000000000000000000000000000"),
	(b"11000001111101100001010001111011", b"11000010101110111101110000101001"), -- -63.17 + -30.76 = -93.93
	(b"11000010101001010101011100001010", b"00000000000000000000000000000000"),
	(b"01000010100001010110101110000101", b"11000001011111110101110000101000"), -- -82.67 + 66.71 = -15.96
	(b"11000010100110101101000111101100", b"00000000000000000000000000000000"),
	(b"00111111101100001010001111010111", b"11000010100110000000111101011101"), -- -77.41 + 1.38 = -76.03
	(b"01000010100000111100011110101110", b"00000000000000000000000000000000"),
	(b"11000001001011010111000010100100", b"01000010010111000011001100110011"), -- 65.89 + -10.84 = 55.05
	(b"11000010011000110101000111101100", b"00000000000000000000000000000000"),
	(b"11000010101111010001010001111011", b"11000011000101110101111010111000"), -- -56.83 + -94.54 = -151.37
	(b"01000010011100100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110111101011100001010001111", b"01000010011100000010100011110110"), -- 60.52 + -0.48 = 60.04
	(b"11000000011000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000111000010100011110110", b"11000000101111111010111000010100"), -- -3.55 + -2.44 = -5.99
	(b"01000010100101100100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001010110001111010111000", b"01000010111010111101110000101001"), -- 75.15 + 42.78 = 117.93
	(b"11000010011110001111010111000011", b"00000000000000000000000000000000"),
	(b"11000010010001001110000101001000", b"11000010110111101110101110000110"), -- -62.24 + -49.22 = -111.46
	(b"11000010001101010111101011100001", b"00000000000000000000000000000000"),
	(b"01000001111111001000111101011100", b"11000001010111001100110011001100"), -- -45.37 + 31.57 = -13.8
	(b"01000001010001001111010111000011", b"00000000000000000000000000000000"),
	(b"11000010001011110000000000000000", b"11000001111110111000010100011110"), -- 12.31 + -43.75 = -31.44
	(b"01000010000001011000111101011100", b"00000000000000000000000000000000"),
	(b"01000001101011011000010100011111", b"01000010010111000101000111101100"), -- 33.39 + 21.69 = 55.08
	(b"01000010101010101000101000111101", b"00000000000000000000000000000000"),
	(b"11000010001000110000000000000000", b"01000010001100100001010001111010"), -- 85.27 + -40.75 = 44.52
	(b"01000010010101101011100001010010", b"00000000000000000000000000000000"),
	(b"01000010010001001100110011001101", b"01000010110011011100001010010000"), -- 53.68 + 49.2 = 102.88
	(b"11000001001110110000101000111101", b"00000000000000000000000000000000"),
	(b"01000010010101001011100001010010", b"01000010001001011111010111000011"), -- -11.69 + 53.18 = 41.49
	(b"01000010000101111110000101001000", b"00000000000000000000000000000000"),
	(b"11000010101001101010111000010100", b"11000010001101010111101011100000"), -- 37.97 + -83.34 = -45.37
	(b"11000010100100101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010011110110111000010100100", b"11000001001010011110101110001000"), -- -73.48 + 62.86 = -10.62
	(b"11000010000000110001111010111000", b"00000000000000000000000000000000"),
	(b"11000010001001110111101011100001", b"11000010100101010100110011001100"), -- -32.78 + -41.87 = -74.65
	(b"01000001000100010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000101101111010111000010100", b"01000000010101100110011001101000"), -- 9.09 + -5.74 = 3.35
	(b"11000010100110001111101011100001", b"00000000000000000000000000000000"),
	(b"01000010100110111010001111010111", b"00111111101010100011110110000000"), -- -76.49 + 77.82 = 1.33
	(b"01000001101101010000101000111101", b"00000000000000000000000000000000"),
	(b"11000001100010100001010001111011", b"01000000101010111101011100001000"), -- 22.63 + -17.26 = 5.37
	(b"11000010101111101011110101110001", b"00000000000000000000000000000000"),
	(b"11000010100011011101011100001010", b"11000011001001100100101000111110"), -- -95.37 + -70.92 = -166.29
	(b"11000010010011110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000001110111000010100100", b"11000010101010110011100001010010"), -- -51.75 + -33.86 = -85.61
	(b"01000001111100000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011011010011001100110011", b"01000010101100101011001100110011"), -- 30.05 + 59.3 = 89.35
	(b"11000001101111010000101000111101", b"00000000000000000000000000000000"),
	(b"11000010000101101110000101001000", b"11000010011101010110011001100110"), -- -23.63 + -37.72 = -61.35
	(b"01000010000111100111000010100100", b"00000000000000000000000000000000"),
	(b"11000010100011011001100110011010", b"11000001111110011000010100100000"), -- 39.61 + -70.8 = -31.19
	(b"01000010101110001010100011110110", b"00000000000000000000000000000000"),
	(b"01000010101001011100001010001111", b"01000011001011110011010111000010"), -- 92.33 + 82.88 = 175.21
	(b"01000001111110100010100011110110", b"00000000000000000000000000000000"),
	(b"01000010110000011000000000000000", b"01000011000000000000010100011111"), -- 31.27 + 96.75 = 128.02
	(b"01000000111011000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"01000000010001011100001010001110"), -- 7.39 + -4.3 = 3.09
	(b"01000010101101110011110101110001", b"00000000000000000000000000000000"),
	(b"01000000101101010111000010100100", b"01000010110000101001010001111011"), -- 91.62 + 5.67 = 97.29
	(b"11000010101110010010001111010111", b"00000000000000000000000000000000"),
	(b"11000010101101110010111000010100", b"11000011001110000010100011110110"), -- -92.57 + -91.59 = -184.16
	(b"11000010001101100010100011110110", b"00000000000000000000000000000000"),
	(b"11000001101100001011100001010010", b"11000010100001110100001010010000"), -- -45.54 + -22.09 = -67.63
	(b"01000010100011000100001010001111", b"00000000000000000000000000000000"),
	(b"11000001100001101000111101011100", b"01000010010101010011110101110000"), -- 70.13 + -16.82 = 53.31
	(b"01000000100101100001010001111011", b"00000000000000000000000000000000"),
	(b"01000001011000101011100001010010", b"01000001100101101110000101001000"), -- 4.69 + 14.17 = 18.86
	(b"11000001100010100010100011110110", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"11000001100001111010111000010101"), -- -17.27 + 0.31 = -16.96
	(b"11000010011010101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001000011111010111000011", b"11000001100100010100011110101110"), -- -58.65 + 40.49 = -18.16
	(b"01000010100000110000111101011100", b"00000000000000000000000000000000"),
	(b"01000010010111100111101011100001", b"01000010111100100100110011001100"), -- 65.53 + 55.62 = 121.15
	(b"01000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000010100010000100011110101110", b"01000010100011110001111010111000"), -- 3.42 + 68.14 = 71.56
	(b"11000001011110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000010101100110110101110000101", b"01000010100101000110000101001000"), -- -15.52 + 89.71 = 74.19
	(b"11000001100010110000101000111101", b"00000000000000000000000000000000"),
	(b"01000010101011001110011001100110", b"01000010100010100010001111010111"), -- -17.38 + 86.45 = 69.07
	(b"01000001111001111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010110001001011110101110001", b"01000010111111101001111010111001"), -- 28.94 + 98.37 = 127.31
	(b"11000010101000011001111010111000", b"00000000000000000000000000000000"),
	(b"01000010011011101100001010001111", b"11000001101010001111010111000010"), -- -80.81 + 59.69 = -21.12
	(b"01000010100000101100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100011011000000000000000", b"01000011000010000010000101001000"), -- 65.38 + 70.75 = 136.13
	(b"01000001011100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101101110101110000101001", b"11000010100110010100001010001111"), -- 15.05 + -91.68 = -76.63
	(b"11000010100011101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010101111101010001111010111", b"01000001101111101011100001010000"), -- -71.48 + 95.32 = 23.84
	(b"01000001001101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000010000110011011100001010010", b"11000001110110010011001100110100"), -- 11.28 + -38.43 = -27.15
	(b"01000010101101011001010001111011", b"00000000000000000000000000000000"),
	(b"01000001100110000001010001111011", b"01000010110110111001100110011010"), -- 90.79 + 19.01 = 109.8
	(b"01000010011010001100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100100011000010100011111", b"01000011000000101111001100110011"), -- 58.19 + 72.76 = 130.95
	(b"01000010101111110111010111000011", b"00000000000000000000000000000000"),
	(b"11000001011111101000111101011100", b"01000010100111111010001111011000"), -- 95.73 + -15.91 = 79.82
	(b"01000010010010110101110000101001", b"00000000000000000000000000000000"),
	(b"11000010101000010110000101001000", b"11000001111011101100110011001110"), -- 50.84 + -80.69 = -29.85
	(b"01000010011001110001111010111000", b"00000000000000000000000000000000"),
	(b"01000010101000100001100110011010", b"01000011000010101101010001111011"), -- 57.78 + 81.05 = 138.83
	(b"01000010011011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101111101011100001010", b"01000010010010010011110101110000"), -- 59.8 + -9.49 = 50.31
	(b"01000001000101101110000101001000", b"00000000000000000000000000000000"),
	(b"11000010010110010000101000111101", b"11000010001100110101000111101011"), -- 9.43 + -54.26 = -44.83
	(b"11000010011110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000010001010110101110000101001", b"11000010110100110111000010100100"), -- -62.88 + -42.84 = -105.72
	(b"01000010100101101110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000011101000010100011111", b"01000010000111110100011110101101"), -- 75.45 + -35.63 = 39.82
	(b"11000001101110011100001010001111", b"00000000000000000000000000000000"),
	(b"01000010101010001101011100001010", b"01000010011101001100110011001100"), -- -23.22 + 84.42 = 61.2
	(b"11000010100001111110000101001000", b"00000000000000000000000000000000"),
	(b"11000000111011000111101011100001", b"11000010100101101010100011110110"), -- -67.94 + -7.39 = -75.33
	(b"01000010101111011001111010111000", b"00000000000000000000000000000000"),
	(b"11000010101111110111000010100100", b"10111111011010001111011000000000"), -- 94.81 + -95.72 = -0.910004
	(b"01000010001100000001010001111011", b"00000000000000000000000000000000"),
	(b"00111111110101000111101011100001", b"01000010001101101011100001010010"), -- 44.02 + 1.66 = 45.68
	(b"11000010110001110001010001111011", b"00000000000000000000000000000000"),
	(b"11000010000001010001010001111011", b"11000011000001001100111101011100"), -- -99.54 + -33.27 = -132.81
	(b"11000010010101001100001010001111", b"00000000000000000000000000000000"),
	(b"11000010001010101101011100001010", b"11000010101111111100110011001100"), -- -53.19 + -42.71 = -95.9
	(b"11000010100001001101000111101100", b"00000000000000000000000000000000"),
	(b"01000010101010000101011100001010", b"01000001100011100001010001111000"), -- -66.41 + 84.17 = 17.76
	(b"01000001110111110000101000111101", b"00000000000000000000000000000000"),
	(b"11000001100011000101000111101100", b"01000001001001010111000010100010"), -- 27.88 + -17.54 = 10.34
	(b"01000010011110010101110000101001", b"00000000000000000000000000000000"),
	(b"11000010010010001111010111000011", b"01000001010000011001100110011000"), -- 62.34 + -50.24 = 12.1
	(b"11000010010011110001010001111011", b"00000000000000000000000000000000"),
	(b"01000010010001010111101011100001", b"11000000000110011001100110100000"), -- -51.77 + 49.37 = -2.4
	(b"11000010110000110100011110101110", b"00000000000000000000000000000000"),
	(b"11000010000001011001100110011010", b"11000011000000110000101000111110"), -- -97.64 + -33.4 = -131.04
	(b"11000010101000100110101110000101", b"00000000000000000000000000000000"),
	(b"11000001100011000010100011110110", b"11000010110001010111010111000010"), -- -81.21 + -17.52 = -98.73
	(b"01000010100000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011111110111000010100100", b"00111111011100001010010000000000"), -- 64.8 + -63.86 = 0.940002
	(b"11000010011101101000010100011111", b"00000000000000000000000000000000"),
	(b"11000001011001000010100011110110", b"11000010100101111100011110101110"), -- -61.63 + -14.26 = -75.89
	(b"11000010001011111010001111010111", b"00000000000000000000000000000000"),
	(b"11000010011010111101011100001010", b"11000010110011011011110101110000"), -- -43.91 + -58.96 = -102.87
	(b"01000010011110111000111101011100", b"00000000000000000000000000000000"),
	(b"01000010011100011110101110000101", b"01000010111101101011110101110000"), -- 62.89 + 60.48 = 123.37
	(b"11000010100101000010001111010111", b"00000000000000000000000000000000"),
	(b"01000000111111100110011001100110", b"11000010100001000011110101110001"), -- -74.07 + 7.95 = -66.12
	(b"11000010100111001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011011011110101110000101", b"11000001100101101000111101011110"), -- -78.3 + 59.48 = -18.82
	(b"11000010001110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001011101000101000111101100", b"11000010011101111111010111000011"), -- -46.72 + -15.27 = -61.99
	(b"11000001110010010100011110101110", b"00000000000000000000000000000000"),
	(b"11000010000011100111101011100001", b"11000010011100110001111010111000"), -- -25.16 + -35.62 = -60.78
	(b"11000010101011010000101000111101", b"00000000000000000000000000000000"),
	(b"01000001111010000000000000000000", b"11000010011001100001010001111010"), -- -86.52 + 29 = -57.52
	(b"11000010100100010110101110000101", b"00000000000000000000000000000000"),
	(b"01000001001000110011001100110011", b"11000010011110100000101000111101"), -- -72.71 + 10.2 = -62.51
	(b"11000010100000111101000111101100", b"00000000000000000000000000000000"),
	(b"11000001111110111110101110000101", b"11000010110000101100110011001101"), -- -65.91 + -31.49 = -97.4
	(b"11000001110111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001110110111101011100001", b"11000010100101001101011100001010"), -- -27.55 + -46.87 = -74.42
	(b"11000010000100011010111000010100", b"00000000000000000000000000000000"),
	(b"11000010101001111011110101110001", b"11000010111100001001010001111011"), -- -36.42 + -83.87 = -120.29
	(b"11000001100000101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001010101000101000111101100", b"11000001111011010000101000111110"), -- -16.36 + -13.27 = -29.63
	(b"11000010011001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001011101000010100011111", b"11000010110010101010100011110110"), -- -57.7 + -43.63 = -101.33
	(b"01000010101111001000010100011111", b"00000000000000000000000000000000"),
	(b"01000010001101101010111000010100", b"01000011000010111110111000010100"), -- 94.26 + 45.67 = 139.93
	(b"01000001010000000010100011110110", b"00000000000000000000000000000000"),
	(b"01000001101100011101011100001010", b"01000010000010001111010111000010"), -- 12.01 + 22.23 = 34.24
	(b"11000010110001000100011110101110", b"00000000000000000000000000000000"),
	(b"11000010010001101000010100011111", b"11000011000100111100010100011111"), -- -98.14 + -49.63 = -147.77
	(b"11000001100011001010001111010111", b"00000000000000000000000000000000"),
	(b"01000010101011100001010001111011", b"01000010100010101110101110000101"), -- -17.58 + 87.04 = 69.46
	(b"11000010101101011000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101000100001100110011010", b"11000001000110110011001100110000"), -- -90.75 + 81.05 = -9.7
	(b"11000001110001110000101000111101", b"00000000000000000000000000000000"),
	(b"01000001110000100110011001100110", b"10111111000101000111101011100000"), -- -24.88 + 24.3 = -0.58
	(b"11000010100010011011110101110001", b"00000000000000000000000000000000"),
	(b"01000010001100100010100011110110", b"11000001110000101010001111011000"), -- -68.87 + 44.54 = -24.33
	(b"01000010010001100100011110101110", b"00000000000000000000000000000000"),
	(b"11000001101110011010111000010100", b"01000001110100101110000101001000"), -- 49.57 + -23.21 = 26.36
	(b"01000010100010101101011100001010", b"00000000000000000000000000000000"),
	(b"11000001101101111000010100011111", b"01000010001110011110101110000100"), -- 69.42 + -22.94 = 46.48
	(b"01000010010100010100011110101110", b"00000000000000000000000000000000"),
	(b"11000010010011110011001100110011", b"00111111000001010001111011000000"), -- 52.32 + -51.8 = 0.52
	(b"11000010000100110010100011110110", b"00000000000000000000000000000000"),
	(b"01000001100110000000000000000000", b"11000001100011100101000111101100"), -- -36.79 + 19 = -17.79
	(b"11000001110110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100100001000101000111101", b"01000010001100110111101011100000"), -- -27.4 + 72.27 = 44.87
	(b"11000000001101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000010101011000000101000111101", b"11000010101100011100001010001111"), -- -2.86 + -86.02 = -88.88
	(b"11000010001101101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100010000101000111101100", b"11000010111000111011100001010010"), -- -45.7 + -68.16 = -113.86
	(b"11000010001101011010111000010100", b"00000000000000000000000000000000"),
	(b"11000010101111011000101000111101", b"11000011000011000011000010100100"), -- -45.42 + -94.77 = -140.19
	(b"01000010100010100111010111000011", b"00000000000000000000000000000000"),
	(b"01000001000111110000101000111101", b"01000010100111100101011100001011"), -- 69.23 + 9.94 = 79.17
	(b"11000010101001011100011110101110", b"00000000000000000000000000000000"),
	(b"01000010011011100111101011100001", b"11000001101110100010100011110110"), -- -82.89 + 59.62 = -23.27
	(b"11000010011011001011100001010010", b"00000000000000000000000000000000"),
	(b"01000000101111111010111000010100", b"11000010010101001100001010010000"), -- -59.18 + 5.99 = -53.19
	(b"11000010110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100000001110011001100110", b"11000010000001001001100110011010"), -- -97.6 + 64.45 = -33.15
	(b"11000010000101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011000001000111101011100", b"11000010101110110100011110101110"), -- -37.5 + -56.14 = -93.64
	(b"01000010011000101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000100011100110011001100110", b"01000010011101001000010100011111"), -- 56.68 + 4.45 = 61.13
	(b"11000010101100101001111010111000", b"00000000000000000000000000000000"),
	(b"01000010101101111000010100011111", b"01000000000111001100110011100000"), -- -89.31 + 91.76 = 2.45
	(b"01000010101101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001011001010001111010111", b"01000010001110110101110000101001"), -- 90 + -43.16 = 46.84
	(b"01000010011000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000001000101101110000101001000", b"01000010001111001101011100001010"), -- 56.64 + -9.43 = 47.21
	(b"01000010110001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101101010001111010111000", b"01000010101110001010111000010100"), -- 98 + -5.66 = 92.34
	(b"01000000011100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000001111100011110101110000101", b"01000010000010000011001100110011"), -- 3.81 + 30.24 = 34.05
	(b"01000000110000100011110101110001", b"00000000000000000000000000000000"),
	(b"11000010011110001101011100001010", b"11000010011000001000111101011100"), -- 6.07 + -62.21 = -56.14
	(b"01000010101010010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000100100101000111101011100", b"01000010101100100111000010100100"), -- 84.64 + 4.58 = 89.22
	(b"01000010101010111011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101011100001100110011010", b"01000011001011001110011001100110"), -- 85.85 + 87.05 = 172.9
	(b"01000000100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001110101101011100001010", b"11000010001001111101011100001010"), -- 4.75 + -46.71 = -41.96
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010101001110110011001100110", b"01000010101010001010100011110101"), -- 0.63 + 83.7 = 84.33
	(b"01000010100000110100001010001111", b"00000000000000000000000000000000"),
	(b"01000010011001110110011001100110", b"01000010111101101111010111000010"), -- 65.63 + 57.85 = 123.48
	(b"11000010110001111001010001111011", b"00000000000000000000000000000000"),
	(b"11000010001000000010100011110110", b"11000011000010111101010001111011"), -- -99.79 + -40.04 = -139.83
	(b"11000010101010111111000010100100", b"00000000000000000000000000000000"),
	(b"11000001110101110001111010111000", b"11000010111000011011100001010010"), -- -85.97 + -26.89 = -112.86
	(b"11000010011111011010111000010100", b"00000000000000000000000000000000"),
	(b"01000010100100001100001010001111", b"01000001000011110101110000101000"), -- -63.42 + 72.38 = 8.96
	(b"01000010101111110001010001111011", b"00000000000000000000000000000000"),
	(b"01000001011001011110101110000101", b"01000010110110111101000111101100"), -- 95.54 + 14.37 = 109.91
	(b"01000010100111111000010100011111", b"00000000000000000000000000000000"),
	(b"11000001000010010001111010111000", b"01000010100011100110000101001000"), -- 79.76 + -8.57 = 71.19
	(b"01000010100110001000101000111101", b"00000000000000000000000000000000"),
	(b"01000010101100100011001100110011", b"01000011001001010101111010111000"), -- 76.27 + 89.1 = 165.37
	(b"11000010101000100001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111101101100110011001101", b"11000010110111111100110011001101"), -- -81.05 + -30.85 = -111.9
	(b"11000010010111110011110101110001", b"00000000000000000000000000000000"),
	(b"01000010100001111001100110011010", b"01000001001111111101011100001100"), -- -55.81 + 67.8 = 11.99
	(b"01000010101000100110000101001000", b"00000000000000000000000000000000"),
	(b"01000010000010010000101000111101", b"01000010111001101110011001100110"), -- 81.19 + 34.26 = 115.45
	(b"11000010000000001111010111000011", b"00000000000000000000000000000000"),
	(b"11000010010010110001111010111000", b"11000010101001100000101000111110"), -- -32.24 + -50.78 = -83.02
	(b"01000000110000011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010100010000011001100110011", b"01000010100101000101000111101011"), -- 6.06 + 68.1 = 74.16
	(b"11000001101010101010001111010111", b"00000000000000000000000000000000"),
	(b"11000010100011100000111101011100", b"11000010101110001011100001010010"), -- -21.33 + -71.03 = -92.36
	(b"11000010100111000111101011100001", b"00000000000000000000000000000000"),
	(b"11000010001110010010100011110110", b"11000010111110010000111101011100"), -- -78.24 + -46.29 = -124.53
	(b"11000010100110111011110101110001", b"00000000000000000000000000000000"),
	(b"01000010001100010000000000000000", b"11000010000001100111101011100010"), -- -77.87 + 44.25 = -33.62
	(b"01000010100101100111000010100100", b"00000000000000000000000000000000"),
	(b"11000001110011100110011001100110", b"01000010010001011010111000010101"), -- 75.22 + -25.8 = 49.42
	(b"11000010011010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000010001010110010100011110110", b"11000001011111101110000101001000"), -- -58.72 + 42.79 = -15.93
	(b"01000010101100100100001010001111", b"00000000000000000000000000000000"),
	(b"01000010101010000101011100001010", b"01000011001011010100110011001100"), -- 89.13 + 84.17 = 173.3
	(b"01000010000101001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010000101111110101110000101", b"01000010100101100011110101110000"), -- 37.14 + 37.98 = 75.12
	(b"11000010001001111100001010001111", b"00000000000000000000000000000000"),
	(b"11000010011101100111000010100100", b"11000010110011110001100110011010"), -- -41.94 + -61.61 = -103.55
	(b"01000010001110100111000010100100", b"00000000000000000000000000000000"),
	(b"01000010011011111101011100001010", b"01000010110101010010001111010111"), -- 46.61 + 59.96 = 106.57
	(b"01000001100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100001011000000000000000", b"11000010010001001001100110011010"), -- 17.6 + -66.75 = -49.15
	(b"11000000101010011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010001001011010001111010111", b"01000010000100000110011001100110"), -- -5.31 + 41.41 = 36.1
	(b"11000010001011010011110101110001", b"00000000000000000000000000000000"),
	(b"01000010101100001111010111000011", b"01000010001101001010111000010101"), -- -43.31 + 88.48 = 45.17
	(b"11000010000100001110000101001000", b"00000000000000000000000000000000"),
	(b"11000001101011001110000101001000", b"11000010011001110101000111101100"), -- -36.22 + -21.61 = -57.83
	(b"01000010100100000100001010001111", b"00000000000000000000000000000000"),
	(b"01000010011010101000010100011111", b"01000011000000101100001010001111"), -- 72.13 + 58.63 = 130.76
	(b"11000010010011010011110101110001", b"00000000000000000000000000000000"),
	(b"11000000101000111000010100011111", b"11000010011000011010111000010101"), -- -51.31 + -5.11 = -56.42
	(b"01000010100000001010100011110110", b"00000000000000000000000000000000"),
	(b"01000010000100010101000111101100", b"01000010110010010101000111101100"), -- 64.33 + 36.33 = 100.66
	(b"01000010011001101100001010001111", b"00000000000000000000000000000000"),
	(b"11000001100001111010111000010100", b"01000010001000101110101110000101"), -- 57.69 + -16.96 = 40.73
	(b"11000001000010001010001111010111", b"00000000000000000000000000000000"),
	(b"11000010001000101110101110000101", b"11000010010001010001010001111011"), -- -8.54 + -40.73 = -49.27
	(b"11000001110100011000010100011111", b"00000000000000000000000000000000"),
	(b"11000010100011001010100011110110", b"11000010110000010000101000111110"), -- -26.19 + -70.33 = -96.52
	(b"01000010110001101000010100011111", b"00000000000000000000000000000000"),
	(b"11000010100100111100110011001101", b"01000001110010101110000101001000"), -- 99.26 + -73.9 = 25.36
	(b"10111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100010110001111010111000", b"11000001100100010001111010111000"), -- -0.75 + -17.39 = -18.14
	(b"01000010011001000101000111101100", b"00000000000000000000000000000000"),
	(b"11000010011110111100110011001101", b"11000000101110111101011100001000"), -- 57.08 + -62.95 = -5.87
	(b"11000010101111001111101011100001", b"00000000000000000000000000000000"),
	(b"11000010110000001011001100110011", b"11000011001111101101011100001010"), -- -94.49 + -96.35 = -190.84
	(b"11000000100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011111100000000000000000", b"11000010100010001000000000000000"), -- -4.75 + -63.5 = -68.25
	(b"11000010100110110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000010101001100011110101110000"), -- -77.52 + -5.6 = -83.12
	(b"01000010001011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001011000111101011100001", b"00111111010001111010111001000000"), -- 43.9 + -43.12 = 0.780003
	(b"11000010110001101111000010100100", b"00000000000000000000000000000000"),
	(b"11000001011001000101000111101100", b"11000010111000110111101011100010"), -- -99.47 + -14.27 = -113.74
	(b"01000010011100010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011100011110101110000101", b"01000010111100011000111101011100"), -- 60.3 + 60.48 = 120.78
	(b"01000010010100101000010100011111", b"00000000000000000000000000000000"),
	(b"11000010100110111001100110011010", b"11000001110010010101110000101010"), -- 52.63 + -77.8 = -25.17
	(b"01000010100101100001111010111000", b"00000000000000000000000000000000"),
	(b"11000010001111111100001010001111", b"01000001110110001111010111000010"), -- 75.06 + -47.94 = 27.12
	(b"01000010011111010100011110101110", b"00000000000000000000000000000000"),
	(b"11000010000110110001010001111011", b"01000001110001000110011001100110"), -- 63.32 + -38.77 = 24.55
	(b"01000010101111010111010111000011", b"00000000000000000000000000000000"),
	(b"11000010100000100000000000000000", b"01000001111011011101011100001100"), -- 94.73 + -65 = 29.73
	(b"11000010101100000110101110000101", b"00000000000000000000000000000000"),
	(b"01000010010010011110000101001000", b"11000010000101101111010111000010"), -- -88.21 + 50.47 = -37.74
	(b"11000010100001101011110101110001", b"00000000000000000000000000000000"),
	(b"11000010100011100000101000111101", b"11000011000010100110001111010111"), -- -67.37 + -71.02 = -138.39
	(b"11000010000101100000101000111101", b"00000000000000000000000000000000"),
	(b"11000010101001100010111000010100", b"11000010111100010011001100110010"), -- -37.51 + -83.09 = -120.6
	(b"01000010011110010000101000111101", b"00000000000000000000000000000000"),
	(b"11000001101111100010100011110110", b"01000010000110011111010111000010"), -- 62.26 + -23.77 = 38.49
	(b"01000010001000010001111010111000", b"00000000000000000000000000000000"),
	(b"01000010100110101011100001010010", b"01000010111010110100011110101110"), -- 40.28 + 77.36 = 117.64
	(b"11000010000001100001111010111000", b"00000000000000000000000000000000"),
	(b"01000010011100101010111000010100", b"01000001110110010001111010111000"), -- -33.53 + 60.67 = 27.14
	(b"11000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111010110011001100110", b"11000010000101101001100110011010"), -- -93 + 55.35 = -37.65
	(b"11000010100100101001100110011010", b"00000000000000000000000000000000"),
	(b"01000001110011001011100001010010", b"11000010001111101101011100001011"), -- -73.3 + 25.59 = -47.71
	(b"11000010010111011111010111000011", b"00000000000000000000000000000000"),
	(b"01000010010001011000111101011100", b"11000000110000110011001100111000"), -- -55.49 + 49.39 = -6.1
	(b"01000001110000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010001111010111000011", b"01000001011101111101011100001001"), -- 24.05 + -8.56 = 15.49
	(b"01000010011000111010001111010111", b"00000000000000000000000000000000"),
	(b"11000010010101110101110000101001", b"01000000010001000111101011100000"), -- 56.91 + -53.84 = 3.07
	(b"01000000111010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100101011110101110000101", b"01000001110011111110101110000101"), -- 7.25 + 18.74 = 25.99
	(b"11000010101001000010001111010111", b"00000000000000000000000000000000"),
	(b"01000010101000011110000101001000", b"10111111100100001010001111000000"), -- -82.07 + 80.94 = -1.13
	(b"11000010000110010111000010100100", b"00000000000000000000000000000000"),
	(b"11000010000101011011100001010010", b"11000010100101111001010001111011"), -- -38.36 + -37.43 = -75.79
	(b"11000010101110111100011110101110", b"00000000000000000000000000000000"),
	(b"01000001101010000110011001100110", b"11000010100100011010111000010100"), -- -93.89 + 21.05 = -72.84
	(b"01000001101010000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001011010000000000000000000", b"01000010000011100011001100110011"), -- 21.05 + 14.5 = 35.55
	(b"01000001001110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011011101010111000010100", b"11000010010000000001010001111010"), -- 11.65 + -59.67 = -48.02
	(b"01000010000110100100011110101110", b"00000000000000000000000000000000"),
	(b"11000010110001010011110101110001", b"11000010011100000011001100110100"), -- 38.57 + -98.62 = -60.05
	(b"01000010001011000010100011110110", b"00000000000000000000000000000000"),
	(b"01000001101001101010001111010111", b"01000010011111110111101011100010"), -- 43.04 + 20.83 = 63.87
	(b"11000010010100010011110101110001", b"00000000000000000000000000000000"),
	(b"11000010101010110011100001010010", b"11000011000010011110101110000101"), -- -52.31 + -85.61 = -137.92
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000001111111011001100110011010", b"11000001111111010111000010100100"), -- 0.02 + -31.7 = -31.68
	(b"11000010001011110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000010101110000101001000", b"11000010000011001010111000010100"), -- -43.85 + 8.68 = -35.17
	(b"11000010001010011011100001010010", b"00000000000000000000000000000000"),
	(b"01000010010001000001111010111000", b"01000000110100110011001100110000"), -- -42.43 + 49.03 = 6.6
	(b"01000010100001010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"01000010100001001110101110000101"), -- 66.64 + -0.18 = 66.46
	(b"01000010001100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101001000011100001010010", b"01000010111111001001111010111000"), -- 44.2 + 82.11 = 126.31
	(b"11000001110001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000000111010111000010100", b"01000001000001101011100001010000"), -- -24.5 + 32.92 = 8.42
	(b"11000010001110100111000010100100", b"00000000000000000000000000000000"),
	(b"11000010010100011100001010001111", b"11000010110001100001100110011010"), -- -46.61 + -52.44 = -99.05
	(b"11000001000001111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010101000101011110101110001", b"01000010100100011100001010010000"), -- -8.49 + 81.37 = 72.88
	(b"11000010100000111011110101110001", b"00000000000000000000000000000000"),
	(b"11000010110001011100110011001101", b"11000011001001001100010100011111"), -- -65.87 + -98.9 = -164.77
	(b"11000010010101010111101011100001", b"00000000000000000000000000000000"),
	(b"11000010011001111010001111010111", b"11000010110111101000111101011100"), -- -53.37 + -57.91 = -111.28
	(b"01000010011011011110000101001000", b"00000000000000000000000000000000"),
	(b"11000001010100001111010111000011", b"01000010001110011010001111010111"), -- 59.47 + -13.06 = 46.41
	(b"11000010000000111000111101011100", b"00000000000000000000000000000000"),
	(b"11000010000010100111101011100001", b"11000010100001110000010100011110"), -- -32.89 + -34.62 = -67.51
	(b"11000010110001100001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110001010000101000111101", b"11000010111101110101110000101001"), -- -99.05 + -24.63 = -123.68
	(b"01000010101100110001111010111000", b"00000000000000000000000000000000"),
	(b"01000001001010110101110000101001", b"01000010110010001000101000111101"), -- 89.56 + 10.71 = 100.27
	(b"01000010101001000100001010001111", b"00000000000000000000000000000000"),
	(b"01000001001100101110000101001000", b"01000010101110101001111010111000"), -- 82.13 + 11.18 = 93.31
	(b"01000010100101110101011100001010", b"00000000000000000000000000000000"),
	(b"01000010101100010110000101001000", b"01000011001001000101110000101001"), -- 75.67 + 88.69 = 164.36
	(b"10111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010011010101011100001010010", b"01000010011001110011001100110011"), -- -0.88 + 58.68 = 57.8
	(b"11000010001110010010100011110110", b"00000000000000000000000000000000"),
	(b"01000001100001100000000000000000", b"11000001111011000101000111101100"), -- -46.29 + 16.75 = -29.54
	(b"01000000111001110101110000101001", b"00000000000000000000000000000000"),
	(b"01000010100011011100001010001111", b"01000010100111000011100001010010"), -- 7.23 + 70.88 = 78.11
	(b"01000010000100000111101011100001", b"00000000000000000000000000000000"),
	(b"01000010101011100010100011110110", b"01000010111101100110011001100110"), -- 36.12 + 87.08 = 123.2
	(b"11000010010100110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001000110000000000000000", b"11000010101110110011001100110011"), -- -52.85 + -40.75 = -93.6
	(b"01000010010110110001010001111011", b"00000000000000000000000000000000"),
	(b"01000010001101000000101000111101", b"01000010110001111000111101011100"), -- 54.77 + 45.01 = 99.78
	(b"01000000110011010001111010111000", b"00000000000000000000000000000000"),
	(b"01000010001010001101011100001010", b"01000010010000100111101011100001"), -- 6.41 + 42.21 = 48.62
	(b"01000010011100111000111101011100", b"00000000000000000000000000000000"),
	(b"11000010100010100111000010100100", b"11000001000001010100011110110000"), -- 60.89 + -69.22 = -8.33
	(b"11000010001011010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000100010000000000000000000", b"11000010000111000100011110101110"), -- -43.32 + 4.25 = -39.07
	(b"11000010100111001000010100011111", b"00000000000000000000000000000000"),
	(b"11000010100011100101110000101001", b"11000011000101010111000010100100"), -- -78.26 + -71.18 = -149.44
	(b"01000001011001110101110000101001", b"00000000000000000000000000000000"),
	(b"11000010110000011011001100110011", b"11000010101001001100011110101110"), -- 14.46 + -96.85 = -82.39
	(b"01000010001101000111000010100100", b"00000000000000000000000000000000"),
	(b"11000001010011010111000010100100", b"01000010000000010001010001111011"), -- 45.11 + -12.84 = 32.27
	(b"11000010101011000011100001010010", b"00000000000000000000000000000000"),
	(b"11000010000000100010100011110110", b"11000010111011010100110011001101"), -- -86.11 + -32.54 = -118.65
	(b"01000010000010110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000010000010001000111101011100"), -- 34.84 + -0.7 = 34.14
	(b"00111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000010011000110001111010111000", b"01000010011010010101110000101001"), -- 1.56 + 56.78 = 58.34
	(b"01000001010100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000011111000111101011100", b"11000001101101011110101110000101"), -- 13.15 + -35.89 = -22.74
	(b"11000010100100001110101110000101", b"00000000000000000000000000000000"),
	(b"11000010100011000101000111101100", b"11000011000011101001111010111000"), -- -72.46 + -70.16 = -142.62
	(b"01000010000000101011100001010010", b"00000000000000000000000000000000"),
	(b"11000010011110111010001111010111", b"11000001111100011101011100001010"), -- 32.68 + -62.91 = -30.23
	(b"01000001011110111010111000010100", b"00000000000000000000000000000000"),
	(b"01000010101010001011001100110011", b"01000010110010000010100011110110"), -- 15.73 + 84.35 = 100.08
	(b"01000010110000010101011100001010", b"00000000000000000000000000000000"),
	(b"01000001101110100101000111101100", b"01000010111011111110101110000101"), -- 96.67 + 23.29 = 119.96
	(b"11000010101000010000111101011100", b"00000000000000000000000000000000"),
	(b"11000001000100001111010111000011", b"11000010101100110010111000010100"), -- -80.53 + -9.06 = -89.59
	(b"01000010110001101100001010001111", b"00000000000000000000000000000000"),
	(b"01000010000100010111000010100100", b"01000011000001111011110101110000"), -- 99.38 + 36.36 = 135.74
	(b"11000001010111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001010110011110101110000101", b"11000001110110110101110000101001"), -- -13.8 + -13.62 = -27.42
	(b"01000000000110100011110101110001", b"00000000000000000000000000000000"),
	(b"11000010010101011011100001010010", b"11000010010011000001010001111011"), -- 2.41 + -53.43 = -51.02
	(b"01000001111111111100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100111001000000000000000", b"01000010110111000111000010100100"), -- 31.97 + 78.25 = 110.22
	(b"11000010000110100100011110101110", b"00000000000000000000000000000000"),
	(b"01000010100100000000010100011111", b"01000010000001011100001010010000"), -- -38.57 + 72.01 = 33.44
	(b"01000001100010111110101110000101", b"00000000000000000000000000000000"),
	(b"01000010101000101001010001111011", b"01000010110001011000111101011100"), -- 17.49 + 81.29 = 98.78
	(b"11000010001001010000101000111101", b"00000000000000000000000000000000"),
	(b"11000010011011000111101011100001", b"11000010110010001100001010001111"), -- -41.26 + -59.12 = -100.38
	(b"01000010010000110101110000101001", b"00000000000000000000000000000000"),
	(b"01000010100011000010100011110110", b"01000010111011011101011100001010"), -- 48.84 + 70.08 = 118.92
	(b"11000010100100010111000010100100", b"00000000000000000000000000000000"),
	(b"01000001000000101011100001010010", b"11000010100000010001100110011010"), -- -72.72 + 8.17 = -64.55
	(b"11000010100100111110000101001000", b"00000000000000000000000000000000"),
	(b"01000010010001000001010001111011", b"11000001110001110101110000101010"), -- -73.94 + 49.02 = -24.92
	(b"11000010100110100010100011110110", b"00000000000000000000000000000000"),
	(b"01000010011110111001100110011010", b"11000001011000101110000101001000"), -- -77.08 + 62.9 = -14.18
	(b"11000010010001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101100101000111101011100", b"11000001110101110000101000111110"), -- -49.2 + 22.32 = -26.88
	(b"11000010100111001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010001100001010001111", b"11000011001000101010111000010100"), -- -78.3 + -84.38 = -162.68
	(b"11000001101111100101000111101100", b"00000000000000000000000000000000"),
	(b"01000010101110100111010111000011", b"01000010100010101110000101001000"), -- -23.79 + 93.23 = 69.44
	(b"01000010100010110100011110101110", b"00000000000000000000000000000000"),
	(b"11000010100000100100011110101110", b"01000000100100000000000000000000"), -- 69.64 + -65.14 = 4.5
	(b"01000010001011011011100001010010", b"00000000000000000000000000000000"),
	(b"11000000001000110011001100110011", b"01000010001000111000010100011111"), -- 43.43 + -2.55 = 40.88
	(b"11000001100111101010001111010111", b"00000000000000000000000000000000"),
	(b"10111111110010111000010100011111", b"11000001101010110101110000101001"), -- -19.83 + -1.59 = -21.42
	(b"01000001100011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001000010100011110110", b"01000010101001111111010111000011"), -- 17.9 + 66.08 = 83.98
	(b"01000001110000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001011011101000111101011100", b"01000010000111000000101000111110"), -- 24.1 + 14.91 = 39.01
	(b"01000010100011001011100001010010", b"00000000000000000000000000000000"),
	(b"11000010100111110000000000000000", b"11000001000100100011110101110000"), -- 70.36 + -79.5 = -9.14
	(b"11000010100001010001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110001010001111010111", b"11000010011001000000101000111110"), -- -66.55 + 9.54 = -57.01
	(b"01000010100110111011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101111111011100001010010", b"01000011001011011011010111000010"), -- 77.85 + 95.86 = 173.71
	(b"01000010100101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110101100101000111101100", b"01000010010001000000101000111110"), -- 75.8 + -26.79 = 49.01
	(b"11000010100011010001010001111011", b"00000000000000000000000000000000"),
	(b"01000010101001010100001010001111", b"01000001010000010111000010100000"), -- -70.54 + 82.63 = 12.09
	(b"11000010100001110111000010100100", b"00000000000000000000000000000000"),
	(b"11000001110110110100011110101110", b"11000010101111100100001010010000"), -- -67.72 + -27.41 = -95.13
	(b"01000010000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000011011100001010001111", b"01000000010101110000101001000000"), -- 38.8 + -35.44 = 3.36
	(b"11000010000101110001111010111000", b"00000000000000000000000000000000"),
	(b"11000001101101011010111000010100", b"11000010011100011111010111000010"), -- -37.78 + -22.71 = -60.49
	(b"11000010010010111111010111000011", b"00000000000000000000000000000000"),
	(b"01000010010110111100110011001101", b"01000000011111010111000010100000"), -- -50.99 + 54.95 = 3.96
	(b"11000000010011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000010100101111111010111000011", b"01000010100100011000010100011111"), -- -3.22 + 75.98 = 72.76
	(b"11000010101001111000101000111101", b"00000000000000000000000000000000"),
	(b"11000010101110010111000010100100", b"11000011001100000111110101110000"), -- -83.77 + -92.72 = -176.49
	(b"11000010011000011011100001010010", b"00000000000000000000000000000000"),
	(b"11000001111111011101011100001010", b"11000010101100000101000111101100"), -- -56.43 + -31.73 = -88.16
	(b"11000000010000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010101100010110101110000101", b"01000010101010110100110011001101"), -- -3.06 + 88.71 = 85.65
	(b"11000010011100101010001111010111", b"00000000000000000000000000000000"),
	(b"01000010100110011010100011110110", b"01000001100000010101110000101010"), -- -60.66 + 76.83 = 16.17
	(b"11000001011011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000010001001011000111101011100", b"01000001110100110111000010100100"), -- -14.96 + 41.39 = 26.43
	(b"01000000111011010111000010100100", b"00000000000000000000000000000000"),
	(b"01000010011001001111010111000011", b"01000010100000010101000111101100"), -- 7.42 + 57.24 = 64.66
	(b"11000010010110001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010101011101010001111010111", b"01000010000001001011100001010010"), -- -54.14 + 87.32 = 33.18
	(b"11000010101001110011100001010010", b"00000000000000000000000000000000"),
	(b"11000010100010000000101000111101", b"11000011000101111010000101001000"), -- -83.61 + -68.02 = -151.63
	(b"01000001001101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101101100011001100110011", b"01000010110011010001100110011001"), -- 11.45 + 91.1 = 102.55
	(b"01000001010000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001010101011001100110011010", b"01000001110010110011001100110100"), -- 12.05 + 13.35 = 25.4
	(b"00111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000001101010110011001100110011", b"11000001101001100101000111101011"), -- 0.61 + -21.4 = -20.79
	(b"11000010101000110001111010111000", b"00000000000000000000000000000000"),
	(b"01000001010011001010001111010111", b"11000010100010011000101000111101"), -- -81.56 + 12.79 = -68.77
	(b"01000010101101000011110101110001", b"00000000000000000000000000000000"),
	(b"01000001110101101100110011001101", b"01000010111010011111000010100100"), -- 90.12 + 26.85 = 116.97
	(b"11000010001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010110000110000000000000000", b"01000010011000100010100011110110"), -- -40.96 + 97.5 = 56.54
	(b"01000001101011001110000101001000", b"00000000000000000000000000000000"),
	(b"01000010011101011000010100011111", b"01000010101001011111101011100010"), -- 21.61 + 61.38 = 82.99
	(b"01000010100001001101011100001010", b"00000000000000000000000000000000"),
	(b"11000010010001110111000010100100", b"01000001100001000111101011100000"), -- 66.42 + -49.86 = 16.56
	(b"11000010000100111100001010001111", b"00000000000000000000000000000000"),
	(b"01000010001110011100001010001111", b"01000001000110000000000000000000"), -- -36.94 + 46.44 = 9.5
	(b"01000010011010010111000010100100", b"00000000000000000000000000000000"),
	(b"11000010110001011011001100110011", b"11000010001000011111010111000010"), -- 58.36 + -98.85 = -40.49
	(b"01000001010101111101011100001010", b"00000000000000000000000000000000"),
	(b"11000010101110101111101011100001", b"11000010101000000000000000000000"), -- 13.49 + -93.49 = -80
	(b"01000001101011010101110000101001", b"00000000000000000000000000000000"),
	(b"11000001110001010100011110101110", b"11000000001111110101110000101000"), -- 21.67 + -24.66 = -2.99
	(b"11000001111100010000101000111101", b"00000000000000000000000000000000"),
	(b"01000010010000010011001100110011", b"01000001100100010101110000101001"), -- -30.13 + 48.3 = 18.17
	(b"11000001001010010111000010100100", b"00000000000000000000000000000000"),
	(b"01000010110000111100110011001101", b"01000010101011101001111010111000"), -- -10.59 + 97.9 = 87.31
	(b"11000010011100011111010111000011", b"00000000000000000000000000000000"),
	(b"11000001110110100010100011110110", b"11000010101011111000010100011111"), -- -60.49 + -27.27 = -87.76
	(b"11000010100101001000010100011111", b"00000000000000000000000000000000"),
	(b"11000010100000011001100110011010", b"11000011000010110000111101011100"), -- -74.26 + -64.8 = -139.06
	(b"11000010001011110001010001111011", b"00000000000000000000000000000000"),
	(b"11000010110000100101011100001010", b"11000011000011001111000010100100"), -- -43.77 + -97.17 = -140.94
	(b"01000001100010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011000100001010001111011", b"01000000010010101110000101000100"), -- 17.3 + -14.13 = 3.17
	(b"01000010100011011001111010111000", b"00000000000000000000000000000000"),
	(b"01000010101110010011110101110001", b"01000011001000110110111000010100"), -- 70.81 + 92.62 = 163.43
	(b"11000001111101000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110100100010100011110110", b"11000010011000110100011110101110"), -- -30.55 + -26.27 = -56.82
	(b"01000001101100100011110101110001", b"00000000000000000000000000000000"),
	(b"11000010000101000100011110101110", b"11000001011011001010001111010110"), -- 22.28 + -37.07 = -14.79
	(b"11000000101011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000111110101110000101001000", b"11000001010101000111101011100010"), -- -5.44 + -7.84 = -13.28
	(b"01000010011011010111000010100100", b"00000000000000000000000000000000"),
	(b"11000010010000111111010111000011", b"01000001001001011110101110000100"), -- 59.36 + -48.99 = 10.37
	(b"01000010011111010000101000111101", b"00000000000000000000000000000000"),
	(b"11000010110001100110000101001000", b"11000010000011111011100001010011"), -- 63.26 + -99.19 = -35.93
	(b"01000001100001011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000011110111000010100011111", b"01000001101001010101110000101001"), -- 16.74 + 3.93 = 20.67
	(b"11000010100011101101110000101001", b"00000000000000000000000000000000"),
	(b"01000010011101110111101011100001", b"11000001000110001111010111000100"), -- -71.43 + 61.87 = -9.56
	(b"01000010100001101000111101011100", b"00000000000000000000000000000000"),
	(b"01000010000011100111000010100100", b"01000010110011011100011110101110"), -- 67.28 + 35.61 = 102.89
	(b"11000010101000110011100001010010", b"00000000000000000000000000000000"),
	(b"11000001100101000010100011110110", b"11000010110010000100001010010000"), -- -81.61 + -18.52 = -100.13
	(b"11000010010011110111101011100001", b"00000000000000000000000000000000"),
	(b"01000010010011111111010111000011", b"00111101111101011100010000000000"), -- -51.87 + 51.99 = 0.120003
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000000100101000111101100", b"01000001111101001010001111011000"), -- -2 + 32.58 = 30.58
	(b"11000010000110110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100110101101011100001010", b"11000010111010000101011100001010"), -- -38.75 + -77.42 = -116.17
	(b"11000010000001101001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001001100110011001101", b"11000010000101110011001100110100"), -- -33.65 + -4.15 = -37.8
	(b"11000001111101111100001010001111", b"00000000000000000000000000000000"),
	(b"01000010001100111011100001010010", b"01000001010111110101110000101010"), -- -30.97 + 44.93 = 13.96
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001000001111010111000011", b"11000010000111101100001010010000"), -- 0.55 + -40.24 = -39.69
	(b"01000010001001001010111000010100", b"00000000000000000000000000000000"),
	(b"11000001110111001110000101001000", b"01000001010110001111010111000000"), -- 41.17 + -27.61 = 13.56
	(b"01000010011100110001111010111000", b"00000000000000000000000000000000"),
	(b"11000001010110001111010111000011", b"01000010001111001110000101000111"), -- 60.78 + -13.56 = 47.22
	(b"11000010101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000001110110011001100110", b"11000010111000111011001100110011"), -- -80 + -33.85 = -113.85
	(b"01000001100100010000101000111101", b"00000000000000000000000000000000"),
	(b"01000010110001110110011001100110", b"01000010111010111010100011110101"), -- 18.13 + 99.7 = 117.83
	(b"01000010101110010001010001111011", b"00000000000000000000000000000000"),
	(b"11000010101010011010001111010111", b"01000000111101110000101001000000"), -- 92.54 + -84.82 = 7.72
	(b"01000010110000100000101000111101", b"00000000000000000000000000000000"),
	(b"11000001110110111110101110000101", b"01000010100010110000111101011100"), -- 97.02 + -27.49 = 69.53
	(b"11000010001100001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010011000100010100011110110", b"01000001010001100110011001101000"), -- -44.14 + 56.54 = 12.4
	(b"01000010101101011010001111010111", b"00000000000000000000000000000000"),
	(b"11000010011110110000101000111101", b"01000001111000000111101011100010"), -- 90.82 + -62.76 = 28.06
	(b"11000010101100111110101110000101", b"00000000000000000000000000000000"),
	(b"01000010010100111010001111010111", b"11000010000101000011001100110011"), -- -89.96 + 52.91 = -37.05
	(b"01000000111010111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010011111101100001010001111", b"01000010100011100001111010111000"), -- 7.37 + 63.69 = 71.06
	(b"01000010101101110100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001101001100001010001111", b"01000010001110011101011100001011"), -- 91.65 + -45.19 = 46.46
	(b"11000010011101100111101011100001", b"00000000000000000000000000000000"),
	(b"01000010000100100101110000101001", b"11000001110010000011110101110000"), -- -61.62 + 36.59 = -25.03
	(b"11000010000000101100001010001111", b"00000000000000000000000000000000"),
	(b"01000010101010001000000000000000", b"01000010010011100011110101110001"), -- -32.69 + 84.25 = 51.56
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011110111010111000010100", b"11000010011001011010111000010100"), -- 5.5 + -62.92 = -57.42
	(b"11000010001011110000101000111101", b"00000000000000000000000000000000"),
	(b"11000010101011111101011100001010", b"11000011000000111010111000010100"), -- -43.76 + -87.92 = -131.68
	(b"01000001001000000010100011110110", b"00000000000000000000000000000000"),
	(b"11000010101000111011110101110001", b"11000010100011111011100001010010"), -- 10.01 + -81.87 = -71.86
	(b"01000010011101111011100001010010", b"00000000000000000000000000000000"),
	(b"11000010110000000111000010100100", b"11000010000010010010100011110110"), -- 61.93 + -96.22 = -34.29
	(b"01000010011100011000111101011100", b"00000000000000000000000000000000"),
	(b"11000010100111111111010111000011", b"11000001100111001011100001010100"), -- 60.39 + -79.98 = -19.59
	(b"11000010110000000000111101011100", b"00000000000000000000000000000000"),
	(b"01000010001101101111010111000011", b"11000010010010010010100011110101"), -- -96.03 + 45.74 = -50.29
	(b"11000010010001101101011100001010", b"00000000000000000000000000000000"),
	(b"01000001111110111100001010001111", b"11000001100100011110101110000101"), -- -49.71 + 31.47 = -18.24
	(b"11000001100101110111000010100100", b"00000000000000000000000000000000"),
	(b"11000010101100111110000101001000", b"11000010110110011011110101110001"), -- -18.93 + -89.94 = -108.87
	(b"01000010010100101110101110000101", b"00000000000000000000000000000000"),
	(b"01000010101111010110000101001000", b"01000011000100110110101110000101"), -- 52.73 + 94.69 = 147.42
	(b"01000010010010110110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110110011110101110000101", b"01000010001100000010100011110101"), -- 50.85 + -6.81 = 44.04
	(b"11000001111010100111101011100001", b"00000000000000000000000000000000"),
	(b"01000000010101100110011001100110", b"11000001110011111010111000010100"), -- -29.31 + 3.35 = -25.96
	(b"01000010100011011111000010100100", b"00000000000000000000000000000000"),
	(b"01000010000110111011100001010010", b"01000010110110111100110011001101"), -- 70.97 + 38.93 = 109.9
	(b"11000010100010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101110110010100011110110", b"01000001110010010111000010100100"), -- -68.4 + 93.58 = 25.18
	(b"11000010100000110011100001010010", b"00000000000000000000000000000000"),
	(b"01000001101110010000101000111101", b"11000010001010011110101110000110"), -- -65.61 + 23.13 = -42.48
	(b"01000010001101110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100010011000101000111101", b"11000001101101110101110000101000"), -- 45.85 + -68.77 = -22.92
	(b"01000010011011011011100001010010", b"00000000000000000000000000000000"),
	(b"01000001111111001110000101001000", b"01000010101101100001010001111011"), -- 59.43 + 31.61 = 91.04
	(b"11000001110100011000010100011111", b"00000000000000000000000000000000"),
	(b"11000000100101110000101000111101", b"11000001111101110100011110101110"), -- -26.19 + -4.72 = -30.91
	(b"01000001001010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101000100101000111101100", b"11000010100011010101000111101100"), -- 10.5 + -81.16 = -70.66
	(b"11000010000010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000010011011110001010001111011", b"11000010101111010100110011001101"), -- -34.88 + -59.77 = -94.65
	(b"01000010000101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000101110111101011100001", b"10111111010111101011100001000000"), -- 37 + -37.87 = -0.869999
	(b"11000001010011011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010100011111100001010001111", b"01000010011011000000101000111101"), -- -12.87 + 71.88 = 59.01
	(b"01000010100000000100011110101110", b"00000000000000000000000000000000"),
	(b"11000010100110111010111000010100", b"11000001010110110011001100110000"), -- 64.14 + -77.84 = -13.7
	(b"11000010101010110111000010100100", b"00000000000000000000000000000000"),
	(b"01000010110001011111000010100100", b"01000001010101000000000000000000"), -- -85.72 + 98.97 = 13.25
	(b"11000001111100111110101110000101", b"00000000000000000000000000000000"),
	(b"01000010101010101010111000010100", b"01000010010110110110011001100110"), -- -30.49 + 85.34 = 54.85
	(b"11000010110000001110000101001000", b"00000000000000000000000000000000"),
	(b"01000010001011010110011001100110", b"11000010010101000101110000101010"), -- -96.44 + 43.35 = -53.09
	(b"11000010010101011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010010001000000000000000000", b"11000000100011110101110000101000"), -- -53.48 + 49 = -4.48
	(b"01000010101011110100110011001101", b"00000000000000000000000000000000"),
	(b"11000001100100010011001100110011", b"01000010100010110000000000000000"), -- 87.65 + -18.15 = 69.5
	(b"01000010101110100100001010001111", b"00000000000000000000000000000000"),
	(b"01000010001011100100011110101110", b"01000011000010001011001100110011"), -- 93.13 + 43.57 = 136.7
	(b"11000001100011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100011001010001111010111", b"01000010010100100111101011100001"), -- -17.7 + 70.32 = 52.62
	(b"01000010000011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111000100000000000000000", b"01000000111001001100110011010000"), -- 35.4 + -28.25 = 7.15
	(b"01000010011001110111000010100100", b"00000000000000000000000000000000"),
	(b"11000001111101101110000101001000", b"01000001110110000000000000000000"), -- 57.86 + -30.86 = 27
	(b"11000010000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011001100010100011110110", b"11000010101111111110000101001000"), -- -38.4 + -57.54 = -95.94
	(b"11000010101011001100011110101110", b"00000000000000000000000000000000"),
	(b"11000010110001101100011110101110", b"11000011001110011100011110101110"), -- -86.39 + -99.39 = -185.78
	(b"11000010010100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010101011110000101001000", b"00111111101111000010100100000000"), -- -52 + 53.47 = 1.47
	(b"01000010011001101001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111000000010100011111", b"11000010000100010111000010100100"), -- 57.65 + -94.01 = -36.36
	(b"11000001110101101000111101011100", b"00000000000000000000000000000000"),
	(b"01000001110001000001010001111011", b"11000000000100111101011100001000"), -- -26.82 + 24.51 = -2.31
	(b"11000010100110111010111000010100", b"00000000000000000000000000000000"),
	(b"01000001100010010100011110101110", b"11000010011100101011100001010001"), -- -77.84 + 17.16 = -60.68
	(b"11000010001011100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111111100001010001111010111", b"11000010001001101011100001010010"), -- -43.56 + 1.88 = -41.68
	(b"01000010101100011001010001111011", b"00000000000000000000000000000000"),
	(b"11000010101110011111010111000011", b"11000000100001100001010010000000"), -- 88.79 + -92.98 = -4.19
	(b"11000001101100010000101000111101", b"00000000000000000000000000000000"),
	(b"01000010101010010101000111101100", b"01000010011110100001111010111010"), -- -22.13 + 84.66 = 62.53
	(b"11000000111011111010111000010100", b"00000000000000000000000000000000"),
	(b"11000010011011100111000010100100", b"11000010100001100011001100110011"), -- -7.49 + -59.61 = -67.1
	(b"01000001101111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000010001111111100001010001111", b"11000001110000010111000010100011"), -- 23.76 + -47.94 = -24.18
	(b"11000010011010110100011110101110", b"00000000000000000000000000000000"),
	(b"01000010101110001000101000111101", b"01000010000001011100110011001100"), -- -58.82 + 92.27 = 33.45
	(b"01000001101100000001010001111011", b"00000000000000000000000000000000"),
	(b"11000010101111001100011110101110", b"11000010100100001100001010001111"), -- 22.01 + -94.39 = -72.38
	(b"11000010011110011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010011101010001010001111011", b"11000010111101111000000000000000"), -- -62.48 + -61.27 = -123.75
	(b"01000001101110000010100011110110", b"00000000000000000000000000000000"),
	(b"11000010100010111100011110101110", b"11000010001110110111101011100001"), -- 23.02 + -69.89 = -46.87
	(b"11000010101000111001111010111000", b"00000000000000000000000000000000"),
	(b"01000010110001100111000010100100", b"01000001100010110100011110110000"), -- -81.81 + 99.22 = 17.41
	(b"01000010011000001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010101010101000010100011111", b"01000011000011010110011001100110"), -- 56.14 + 85.26 = 141.4
	(b"11000001100110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101111110010001111010111", b"11000010111001010011110101110000"), -- -19.05 + -95.57 = -114.62
	(b"11000010100010000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001110100011110101110", b"10111110111010111000010100000000"), -- -68.1 + 67.64 = -0.459999
	(b"11000000110101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110100101110000101001000", b"10111101011101011100001010000000"), -- -6.65 + 6.59 = -0.0599999
	(b"01000010010100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100000010100011110101110", b"01000010100010010001111010111000"), -- 52.4 + 16.16 = 68.56
	(b"01000010101111010111101011100001", b"00000000000000000000000000000000"),
	(b"01000001010000100110011001100110", b"01000010110101011100011110101110"), -- 94.74 + 12.15 = 106.89
	(b"01000010100101001001010001111011", b"00000000000000000000000000000000"),
	(b"01000001001101000000000000000000", b"01000010101010110001010001111011"), -- 74.29 + 11.25 = 85.54
	(b"01000010101010001010100011110110", b"00000000000000000000000000000000"),
	(b"01000010011111111010001111010111", b"01000011000101000011110101110001"), -- 84.33 + 63.91 = 148.24
	(b"11000001100001001000111101011100", b"00000000000000000000000000000000"),
	(b"11000010001100101010111000010100", b"11000010011101001111010111000010"), -- -16.57 + -44.67 = -61.24
	(b"01000010101010010111101011100001", b"00000000000000000000000000000000"),
	(b"11000010110001110001100110011010", b"11000001011011001111010111001000"), -- 84.74 + -99.55 = -14.81
	(b"01000010100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100101001110011001100110", b"00111111110001100110011010000000"), -- 76 + -74.45 = 1.55
	(b"11000010000100010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001010111010100011110101110", b"11000001101100110101110000101001"), -- -36.25 + 13.83 = -22.42
	(b"11000010000011100101000111101100", b"00000000000000000000000000000000"),
	(b"11000010000001010111000010100100", b"11000010100010011110000101001000"), -- -35.58 + -33.36 = -68.94
	(b"11000010100000001101000111101100", b"00000000000000000000000000000000"),
	(b"01000001010100101110000101001000", b"11000010010011001110101110000110"), -- -64.41 + 13.18 = -51.23
	(b"01000010010111011101011100001010", b"00000000000000000000000000000000"),
	(b"01000010010000011010001111010111", b"01000010110011111011110101110000"), -- 55.46 + 48.41 = 103.87
	(b"01000010010011000001111010111000", b"00000000000000000000000000000000"),
	(b"01000001110011011100001010001111", b"01000010100110011000000000000000"), -- 51.03 + 25.72 = 76.75
	(b"11000010010010000111000010100100", b"00000000000000000000000000000000"),
	(b"01000010011101010011110101110001", b"01000001001100110011001100110100"), -- -50.11 + 61.31 = 11.2
	(b"01000001010001111000010100011111", b"00000000000000000000000000000000"),
	(b"01000010100001100011001100110011", b"01000010100111110010001111010111"), -- 12.47 + 67.1 = 79.57
	(b"01000010011111101000111101011100", b"00000000000000000000000000000000"),
	(b"01000001111110000111101011100001", b"01000010101111010110011001100110"), -- 63.64 + 31.06 = 94.7
	(b"11000010101100100111010111000011", b"00000000000000000000000000000000"),
	(b"11000010100000000000010100011111", b"11000011000110010011110101110001"), -- -89.23 + -64.01 = -153.24
	(b"11000010001010000111000010100100", b"00000000000000000000000000000000"),
	(b"01000010011101110101000111101100", b"01000001100111011100001010010000"), -- -42.11 + 61.83 = 19.72
	(b"11000010000101001010111000010100", b"00000000000000000000000000000000"),
	(b"11000010100001111110011001100110", b"11000010110100100011110101110000"), -- -37.17 + -67.95 = -105.12
	(b"11000010101111110011100001010010", b"00000000000000000000000000000000"),
	(b"11000000111100000101000111101100", b"11000010110011100011110101110001"), -- -95.61 + -7.51 = -103.12
	(b"11000010110000001011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101011010101000111101100", b"11000001000110110000101000111000"), -- -96.35 + 86.66 = -9.68999
	(b"11000001001001110000101000111101", b"00000000000000000000000000000000"),
	(b"01000001101101110001111010111000", b"01000001010001110011001100110011"), -- -10.44 + 22.89 = 12.45
	(b"01000010010111111100001010001111", b"00000000000000000000000000000000"),
	(b"11000001010000010111000010100100", b"01000010001011110110011001100110"), -- 55.94 + -12.09 = 43.85
	(b"11000010001111010000101000111101", b"00000000000000000000000000000000"),
	(b"01000010001111001110101110000101", b"10111100111101011100000000000000"), -- -47.26 + 47.23 = -0.0299988
	(b"01000010000011111110101110000101", b"00000000000000000000000000000000"),
	(b"11000000001010101110000101001000", b"01000010000001010011110101110000"), -- 35.98 + -2.67 = 33.31
	(b"11000010101100111100011110101110", b"00000000000000000000000000000000"),
	(b"01000010010011101000010100011111", b"11000010000110010000101000111101"), -- -89.89 + 51.63 = -38.26
	(b"10111111110010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000010011010110111000010100100", b"01000010011001010010100011110110"), -- -1.57 + 58.86 = 57.29
	(b"11000010101101001000101000111101", b"00000000000000000000000000000000"),
	(b"11000001001011100011110101110001", b"11000010110010100101000111101011"), -- -90.27 + -10.89 = -101.16
	(b"11000001111111001110000101001000", b"00000000000000000000000000000000"),
	(b"11000010000100010111000010100100", b"11000010100001111111000010100100"), -- -31.61 + -36.36 = -67.97
	(b"11000001111111001000111101011100", b"00000000000000000000000000000000"),
	(b"01000001111011000101000111101100", b"11000000000000011110101110000000"), -- -31.57 + 29.54 = -2.03
	(b"01000010100010110110101110000101", b"00000000000000000000000000000000"),
	(b"11000010010100001110000101001000", b"01000001100010111110101110000100"), -- 69.71 + -52.22 = 17.49
	(b"11000001110011000101000111101100", b"00000000000000000000000000000000"),
	(b"11000010001110101010111000010100", b"11000010100100000110101110000101"), -- -25.54 + -46.67 = -72.21
	(b"11000010011001110111101011100001", b"00000000000000000000000000000000"),
	(b"01000001111110010011001100110011", b"11000001110101011100001010001111"), -- -57.87 + 31.15 = -26.72
	(b"01000010000110110001111010111000", b"00000000000000000000000000000000"),
	(b"11000010010101001001100110011010", b"11000001011001011110101110001000"), -- 38.78 + -53.15 = -14.37
	(b"01000010101001101010111000010100", b"00000000000000000000000000000000"),
	(b"01000001101100001000111101011100", b"01000010110100101101000111101011"), -- 83.34 + 22.07 = 105.41
	(b"01000010001010110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110001101011100001010010", b"01000010100001110110000101001000"), -- 42.85 + 24.84 = 67.69
	(b"11000010101011110011110101110001", b"00000000000000000000000000000000"),
	(b"01000010101110000000000000000000", b"01000000100011000010100011110000"), -- -87.62 + 92 = 4.38
	(b"11000001001010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000010010101101110000101001000", b"01000010001011000010100011110110"), -- -10.68 + 53.72 = 43.04
	(b"11000010010110111100001010001111", b"00000000000000000000000000000000"),
	(b"01000001111110110100011110101110", b"11000001101111000011110101110000"), -- -54.94 + 31.41 = -23.53
	(b"01000010100110010100001010001111", b"00000000000000000000000000000000"),
	(b"01000010100100111110011001100110", b"01000011000101101001010001111010"), -- 76.63 + 73.95 = 150.58
	(b"11000010101111000010111000010100", b"00000000000000000000000000000000"),
	(b"11000010110001000001111010111000", b"11000011010000000010011001100110"), -- -94.09 + -98.06 = -192.15
	(b"01000010001101010011110101110001", b"00000000000000000000000000000000"),
	(b"01000001111010001111010111000011", b"01000010100101001101110000101001"), -- 45.31 + 29.12 = 74.43
	(b"11000010100100010100011110101110", b"00000000000000000000000000000000"),
	(b"11000001011000010111000010100100", b"11000010101011010111010111000010"), -- -72.64 + -14.09 = -86.73
	(b"11000010000110110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101111100010001111010111", b"01000010011000001110000101001000"), -- -38.85 + 95.07 = 56.22
	(b"11000010001010001010001111010111", b"00000000000000000000000000000000"),
	(b"01000010101000000110000101001000", b"01000010000110000001111010111001"), -- -42.16 + 80.19 = 38.03
	(b"11000001011100111101011100001010", b"00000000000000000000000000000000"),
	(b"11000010100001000111000010100100", b"11000010101000101110101110000101"), -- -15.24 + -66.22 = -81.46
	(b"01000010000000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000001110010110100011110101110", b"01000010011010010111101011100001"), -- 32.96 + 25.41 = 58.37
	(b"01000010011011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100111011001100110011010", b"11000001100110000000000000000010"), -- 59.8 + -78.8 = -19
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000110101000010100011110110", b"11000000110010000101000111101100"), -- 0.37 + -6.63 = -6.26
	(b"01000010001101000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101110101100110011001101", b"01000011000010100111001100110011"), -- 45.05 + 93.4 = 138.45
	(b"11000010100111011001010001111011", b"00000000000000000000000000000000"),
	(b"01000010100001010000101000111101", b"11000001010001000101000111110000"), -- -78.79 + 66.52 = -12.27
	(b"01000010101100000100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000010100011110101110", b"01000000111100000101000111110000"), -- 88.15 + -80.64 = 7.51
	(b"11000010000010001100001010001111", b"00000000000000000000000000000000"),
	(b"11000010000110010000101000111101", b"11000010100100001110011001100110"), -- -34.19 + -38.26 = -72.45
	(b"01000010101101110001111010111000", b"00000000000000000000000000000000"),
	(b"11000010011011000111000010100100", b"01000010000000011100110011001100"), -- 91.56 + -59.11 = 32.45
	(b"11000010100110011100001010001111", b"00000000000000000000000000000000"),
	(b"01000010001001010101000111101100", b"11000010000011100011001100110010"), -- -76.88 + 41.33 = -35.55
	(b"11000001101100110000101000111101", b"00000000000000000000000000000000"),
	(b"01000001010010000101000111101100", b"11000001000111011100001010001110"), -- -22.38 + 12.52 = -9.86
	(b"01000010100010110110101110000101", b"00000000000000000000000000000000"),
	(b"01000001101011000110011001100110", b"01000010101101101000010100011110"), -- 69.71 + 21.55 = 91.26
	(b"01000010101110000110000101001000", b"00000000000000000000000000000000"),
	(b"01000010001101010000000000000000", b"01000011000010010111000010100100"), -- 92.19 + 45.25 = 137.44
	(b"01000010100100000010111000010100", b"00000000000000000000000000000000"),
	(b"11000010101111101111000010100100", b"11000001101110110000101001000000"), -- 72.09 + -95.47 = -23.38
	(b"11000010011011100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001110001110000101001000", b"11000001010101010100011110101100"), -- -59.55 + 46.22 = -13.33
	(b"01000010100101111000111101011100", b"00000000000000000000000000000000"),
	(b"11000010001101100001111010111000", b"01000001111100100000000000000000"), -- 75.78 + -45.53 = 30.25
	(b"01000010101101100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000111001011100001010001111", b"01000010101001111011100001010010"), -- 91.04 + -7.18 = 83.86
	(b"11000010100010001111101011100001", b"00000000000000000000000000000000"),
	(b"11000010010100011110101110000101", b"11000010111100011111000010100100"), -- -68.49 + -52.48 = -120.97
	(b"11000010001100110100011110101110", b"00000000000000000000000000000000"),
	(b"11000010101001000011100001010010", b"11000010111111011101110000101001"), -- -44.82 + -82.11 = -126.93
	(b"11000010011100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010110000100000010100011111", b"01000010000100100000101000111110"), -- -60.5 + 97.01 = 36.51
	(b"01000010100110110010111000010100", b"00000000000000000000000000000000"),
	(b"11000001010000111101011100001010", b"01000010100000101011001100110011"), -- 77.59 + -12.24 = 65.35
	(b"01000001111010010111000010100100", b"00000000000000000000000000000000"),
	(b"11000010100011101111101011100001", b"11000010001010010011110101110000"), -- 29.18 + -71.49 = -42.31
	(b"01000010101101101001010001111011", b"00000000000000000000000000000000"),
	(b"11000010001011101011100001010010", b"01000010001111100111000010100100"), -- 91.29 + -43.68 = 47.61
	(b"01000010100011000100011110101110", b"00000000000000000000000000000000"),
	(b"11000010011011000111101011100001", b"01000001001100000101000111101100"), -- 70.14 + -59.12 = 11.02
	(b"01000010100010010101000111101100", b"00000000000000000000000000000000"),
	(b"11000010001000000110011001100110", b"01000001111001000111101011100100"), -- 68.66 + -40.1 = 28.56
	(b"11000010010011101110101110000101", b"00000000000000000000000000000000"),
	(b"11000010011001011001100110011010", b"11000010110110100100001010010000"), -- -51.73 + -57.4 = -109.13
	(b"01000001101110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000010101001001001100110011010", b"01000010110100110101000111101100"), -- 23.36 + 82.3 = 105.66
	(b"11000010101001101010001111010111", b"00000000000000000000000000000000"),
	(b"01000001010111001100110011001101", b"11000010100010110000101000111101"), -- -83.32 + 13.8 = -69.52
	(b"01000010001010000001010001111011", b"00000000000000000000000000000000"),
	(b"01000010101010111100110011001101", b"01000010111111111101011100001010"), -- 42.02 + 85.9 = 127.92
	(b"01000010100001011000101000111101", b"00000000000000000000000000000000"),
	(b"11000010101011111000000000000000", b"11000001101001111101011100001100"), -- 66.77 + -87.75 = -20.98
	(b"01000010101011010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100110101010001111010111", b"01000001000100101110000101001000"), -- 86.5 + -77.32 = 9.18
	(b"01000010011011101100001010001111", b"00000000000000000000000000000000"),
	(b"11000010101010110100110011001101", b"11000001110011111010111000010110"), -- 59.69 + -85.65 = -25.96
	(b"01000010101011100101011100001010", b"00000000000000000000000000000000"),
	(b"11000010100011100000101000111101", b"01000001100000010011001100110100"), -- 87.17 + -71.02 = 16.15
	(b"01000001100111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000001111101011110101110000101", b"11000001001011111010111000010100"), -- 19.76 + -30.74 = -10.98
	(b"11000001111111011000010100011111", b"00000000000000000000000000000000"),
	(b"11000010011010101000111101011100", b"11000010101101001010100011110110"), -- -31.69 + -58.64 = -90.33
	(b"11000001100101001011100001010010", b"00000000000000000000000000000000"),
	(b"11000010000010101101011100001010", b"11000010010101010011001100110011"), -- -18.59 + -34.71 = -53.3
	(b"11000010100010010001010001111011", b"00000000000000000000000000000000"),
	(b"11000010110000110000000000000000", b"11000011001001100000101000111110"), -- -68.54 + -97.5 = -166.04
	(b"11000010100011010101110000101001", b"00000000000000000000000000000000"),
	(b"11000001100000001010001111010111", b"11000010101011011000010100011111"), -- -70.68 + -16.08 = -86.76
	(b"01000000101100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000010001010100001010001111011", b"11000010000101000000000000000000"), -- 5.52 + -42.52 = -37
	(b"01000010100000000001111010111000", b"00000000000000000000000000000000"),
	(b"11000010100000101111000010100100", b"10111111101101000111101100000000"), -- 64.06 + -65.47 = -1.41
	(b"01000010100100010011110101110001", b"00000000000000000000000000000000"),
	(b"01000010100110000011100001010010", b"01000011000101001011101011100010"), -- 72.62 + 76.11 = 148.73
	(b"01000010101011010001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000000100111000010100100", b"01000010010101111100001010010000"), -- 86.55 + -32.61 = 53.94
	(b"01000001101111100111101011100001", b"00000000000000000000000000000000"),
	(b"11000010010011000001010001111011", b"11000001110110011010111000010101"), -- 23.81 + -51.02 = -27.21
	(b"01000010110001011111101011100001", b"00000000000000000000000000000000"),
	(b"01000010001001110101000111101100", b"01000011000011001101000111101100"), -- 98.99 + 41.83 = 140.82
	(b"01000010000001110000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110011110101110000101001", b"01000001110110100010100011110110"), -- 33.75 + -6.48 = 27.27
	(b"11000010100110101110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000011001100110011001101", b"11000010111000010100110011001100"), -- -77.45 + -35.2 = -112.65
	(b"01000010001110110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000110001010001111010111000", b"01000010001000100110011001100110"), -- 46.76 + -6.16 = 40.6
	(b"11000010101001110010100011110110", b"00000000000000000000000000000000"),
	(b"01000010001101100101110000101001", b"11000010000101111111010111000011"), -- -83.58 + 45.59 = -37.99
	(b"11000010101111010010100011110110", b"00000000000000000000000000000000"),
	(b"11000010101101101010100011110110", b"11000011001110011110100011110110"), -- -94.58 + -91.33 = -185.91
	(b"01000010010111001011100001010010", b"00000000000000000000000000000000"),
	(b"01000001101000111110101110000101", b"01000010100101110101011100001010"), -- 55.18 + 20.49 = 75.67
	(b"11000010101101111001010001111011", b"00000000000000000000000000000000"),
	(b"01000010110000000100011110101110", b"01000000100010110011001100110000"), -- -91.79 + 96.14 = 4.35
	(b"11000010100001110011100001010010", b"00000000000000000000000000000000"),
	(b"01000010011011100011110101110001", b"11000001000000001100110011001100"), -- -67.61 + 59.56 = -8.05
	(b"01000010101110000110000101001000", b"00000000000000000000000000000000"),
	(b"11000010010001111011100001010010", b"01000010001010010000101000111110"), -- 92.19 + -49.93 = 42.26
	(b"01000010010110100010100011110110", b"00000000000000000000000000000000"),
	(b"01000001011100111010111000010100", b"01000010100010111000101000111110"), -- 54.54 + 15.23 = 69.77
	(b"11000001100110001000111101011100", b"00000000000000000000000000000000"),
	(b"01000010010111101111010111000011", b"01000010000100101010111000010101"), -- -19.07 + 55.74 = 36.67
	(b"11000010001101010001010001111011", b"00000000000000000000000000000000"),
	(b"11000010101010000100110011001101", b"11000011000000010110101110000101"), -- -45.27 + -84.15 = -129.42
	(b"01000010010000111010111000010100", b"00000000000000000000000000000000"),
	(b"11000010000110101111010111000011", b"01000001001000101110000101000100"), -- 48.92 + -38.74 = 10.18
	(b"01000001001000011100001010001111", b"00000000000000000000000000000000"),
	(b"01000010000110110101110000101001", b"01000010010000111100110011001101"), -- 10.11 + 38.84 = 48.95
	(b"01000010001010000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011011001111010111000011", b"01000001110110100101000111101010"), -- 42.1 + -14.81 = 27.29
	(b"11000010101101110111000010100100", b"00000000000000000000000000000000"),
	(b"01000010010011101000010100011111", b"11000010001000000101110000101001"), -- -91.72 + 51.63 = -40.09
	(b"11000001101100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011110111000010100100", b"11000010110111000000101000111110"), -- -22.3 + -87.72 = -110.02
	(b"01000010010001110100011110101110", b"00000000000000000000000000000000"),
	(b"11000001111101000010100011110110", b"01000001100110100110011001100110"), -- 49.82 + -30.52 = 19.3
	(b"11000000110010010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010101110110001100110011010", b"01000010101011101000010100011111"), -- -6.29 + 93.55 = 87.26
	(b"11000010011101011110101110000101", b"00000000000000000000000000000000"),
	(b"11000001111011010101110000101001", b"11000010101101100100110011001101"), -- -61.48 + -29.67 = -91.15
	(b"11000010110000110110101110000101", b"00000000000000000000000000000000"),
	(b"01000010001001100011110101110001", b"11000010011000001001100110011001"), -- -97.71 + 41.56 = -56.15
	(b"01000010101000100110101110000101", b"00000000000000000000000000000000"),
	(b"01000000001011101011100001010010", b"01000010101001111110000101001000"), -- 81.21 + 2.73 = 83.94
	(b"11000000100100000101000111101100", b"00000000000000000000000000000000"),
	(b"01000010000101001100110011001101", b"01000010000000101100001010010000"), -- -4.51 + 37.2 = 32.69
	(b"11000010100111101111000010100100", b"00000000000000000000000000000000"),
	(b"01000010110000000000101000111101", b"01000001100001000110011001100100"), -- -79.47 + 96.02 = 16.55
	(b"01000001100110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000001101110100110011001100110", b"01000010001010010101110000101001"), -- 19.04 + 23.3 = 42.34
	(b"01000001110110100001010001111011", b"00000000000000000000000000000000"),
	(b"01000010101000100101110000101001", b"01000010110110001110000101001000"), -- 27.26 + 81.18 = 108.44
	(b"01000010101101011000101000111101", b"00000000000000000000000000000000"),
	(b"11000010010100011110101110000101", b"01000010000110010010100011110101"), -- 90.77 + -52.48 = 38.29
	(b"11000010100110111111101011100001", b"00000000000000000000000000000000"),
	(b"11000010100110111001111010111000", b"11000011000110111100110011001100"), -- -77.99 + -77.81 = -155.8
	(b"11000010100100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100011111101011100001010", b"11000011000100000101000111101100"), -- -72.4 + -71.92 = -144.32
	(b"01000010100000000010100011110110", b"00000000000000000000000000000000"),
	(b"01000001101110000010100011110110", b"01000010101011100011001100110100"), -- 64.08 + 23.02 = 87.1
	(b"01000001111111011101011100001010", b"00000000000000000000000000000000"),
	(b"01000001001111011001100110011010", b"01000010001011100101000111101100"), -- 31.73 + 11.85 = 43.58
	(b"01000001111010011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010001111101100110011001101", b"11000001100100111010111000010101"), -- 29.24 + -47.7 = -18.46
	(b"01000010101001011111010111000011", b"00000000000000000000000000000000"),
	(b"11000010110000001000010100011111", b"11000001010101000111101011100000"), -- 82.98 + -96.26 = -13.28
	(b"11000000001001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000010000101011111010111000011", b"01000010000010110111101011100010"), -- -2.62 + 37.49 = 34.87
	(b"01000010101110110001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010111010001111010111", b"01000011001100110101111010111000"), -- 93.55 + 85.82 = 179.37
	(b"01000001110101100010100011110110", b"00000000000000000000000000000000"),
	(b"11000001101101001111010111000011", b"01000000100001001100110011001100"), -- 26.77 + -22.62 = 4.15
	(b"01000010101101101111101011100001", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"01000010101101101011001100110011"), -- 91.49 + -0.14 = 91.35
	(b"01000010100000010001111010111000", b"00000000000000000000000000000000"),
	(b"01000010000101010011001100110011", b"01000010110010111011100001010010"), -- 64.56 + 37.3 = 101.86
	(b"01000000000001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000010101001001101000111101100", b"01000010101010001111101011100010"), -- 2.08 + 82.41 = 84.49
	(b"11000001101100000101000111101100", b"00000000000000000000000000000000"),
	(b"01000010100100011110011001100110", b"01000010010010111010001111010110"), -- -22.04 + 72.95 = 50.91
	(b"01000010100000111010001111010111", b"00000000000000000000000000000000"),
	(b"01000001110111010011001100110011", b"01000010101110101111000010100100"), -- 65.82 + 27.65 = 93.47
	(b"01000001110011010001111010111000", b"00000000000000000000000000000000"),
	(b"01000010100001001010111000010100", b"01000010101101111111010111000010"), -- 25.64 + 66.34 = 91.98
	(b"11000010000101010100011110101110", b"00000000000000000000000000000000"),
	(b"11000001111011001100110011001101", b"11000010100001011101011100001010"), -- -37.32 + -29.6 = -66.92
	(b"01000010101100011001111010111000", b"00000000000000000000000000000000"),
	(b"01000010000000001001100110011010", b"01000010111100011110101110000101"), -- 88.81 + 32.15 = 120.96
	(b"01000010010001000001010001111011", b"00000000000000000000000000000000"),
	(b"11000001011010011100001010001111", b"01000010000010011010001111010111"), -- 49.02 + -14.61 = 34.41
	(b"11000010001000110111101011100001", b"00000000000000000000000000000000"),
	(b"01000001010101000000000000000000", b"11000001110111001111010111000010"), -- -40.87 + 13.25 = -27.62
	(b"11000010000011110010100011110110", b"00000000000000000000000000000000"),
	(b"01000001110000001000111101011100", b"11000001001110111000010100100000"), -- -35.79 + 24.07 = -11.72
	(b"11000001011111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010110000101110000101001", b"11000010100010111010111000010100"), -- -15.75 + -54.09 = -69.84
	(b"01000001011111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110001111001100110011010", b"11000001000100000000000000000001"), -- 15.95 + -24.95 = -9
	(b"01000010101110000101011100001010", b"00000000000000000000000000000000"),
	(b"11000001100110101000111101011100", b"01000010100100011011001100110011"), -- 92.17 + -19.32 = 72.85
	(b"01000000011101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000010011111110010100011110110", b"11000010011011111100110011001101"), -- 3.84 + -63.79 = -59.95
	(b"01000010100100000001111010111000", b"00000000000000000000000000000000"),
	(b"11000000000100101000111101011100", b"01000010100010111000101000111101"), -- 72.06 + -2.29 = 69.77
	(b"11000010100000111000101000111101", b"00000000000000000000000000000000"),
	(b"11000010100011011001010001111011", b"11000011000010001000111101011100"), -- -65.77 + -70.79 = -136.56
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110011111010111000011", b"11000010100011110010100011110110"), -- 5.4 + -76.98 = -71.58
	(b"01000010000010110110011001100110", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"01000010000010011010001111010111"), -- 34.85 + -0.44 = 34.41
	(b"01000001110111000001010001111011", b"00000000000000000000000000000000"),
	(b"01000010000111011100110011001101", b"01000010100001011110101110000101"), -- 27.51 + 39.45 = 66.96
	(b"01000010100100110000010100011111", b"00000000000000000000000000000000"),
	(b"11000001101101000000000000000000", b"01000010010011000000101000111110"), -- 73.51 + -22.5 = 51.01
	(b"01000010011010111110101110000101", b"00000000000000000000000000000000"),
	(b"11000010001101010000101000111101", b"01000001010110111000010100100000"), -- 58.98 + -45.26 = 13.72
	(b"11000010110001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010011001000010100011111", b"11000011000101010101010001111011"), -- -98.2 + -51.13 = -149.33
	(b"11000000110100010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010001000101100001010001111", b"01000010000010001001100110011001"), -- -6.54 + 40.69 = 34.15
	(b"11000010101001011010001111010111", b"00000000000000000000000000000000"),
	(b"01000001011010101110000101001000", b"11000010100010000100011110101110"), -- -82.82 + 14.68 = -68.14
	(b"01000001111011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000010100111000111000010100100", b"11000010010000010011001100110100"), -- 29.92 + -78.22 = -48.3
	(b"01000010100000111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101100110010111000010100", b"01000011000110110111110101110000"), -- 65.9 + 89.59 = 155.49
	(b"01000001101111011101011100001010", b"00000000000000000000000000000000"),
	(b"01000010010110110001111010111000", b"01000010100111010000010100011110"), -- 23.73 + 54.78 = 78.51
	(b"11000001111101010111000010100100", b"00000000000000000000000000000000"),
	(b"01000010100011110000111101011100", b"01000010001000110110011001100110"), -- -30.68 + 71.53 = 40.85
	(b"11000010010101011000010100011111", b"00000000000000000000000000000000"),
	(b"01000010010001100111101011100001", b"11000000011100001010001111100000"), -- -53.38 + 49.62 = -3.76
	(b"01000010000000110101110000101001", b"00000000000000000000000000000000"),
	(b"11000001001101101110000101001000", b"01000001101010110100011110101110"), -- 32.84 + -11.43 = 21.41
	(b"01000010110001111001111010111000", b"00000000000000000000000000000000"),
	(b"11000010100001100110000101001000", b"01000010000000100111101011100000"), -- 99.81 + -67.19 = 32.62
	(b"11000010100101110101011100001010", b"00000000000000000000000000000000"),
	(b"11000010000000010001111010111000", b"11000010110101111110011001100110"), -- -75.67 + -32.28 = -107.95
	(b"01000010011110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000110001111010111000011", b"01000001101111100001010001111010"), -- 62 + -38.24 = 23.76
	(b"11000000101000100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000111001011100001010001111", b"01000000000001110000101000111100"), -- -5.07 + 7.18 = 2.11
	(b"11000010100010100111101011100001", b"00000000000000000000000000000000"),
	(b"11000010101011111111000010100100", b"11000011000111010011010111000010"), -- -69.24 + -87.97 = -157.21
	(b"01000010011110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011000100101000111101100", b"01000000110010100011110101110000"), -- 62.9 + -56.58 = 6.32
	(b"11000010101000101110101110000101", b"00000000000000000000000000000000"),
	(b"01000001101010011000010100011111", b"11000010011100010001010001111010"), -- -81.46 + 21.19 = -60.27
	(b"11000010011000110111000010100100", b"00000000000000000000000000000000"),
	(b"11000010101011100001111010111000", b"11000011000011111110101110000101"), -- -56.86 + -87.06 = -143.92
	(b"11000010010001011000010100011111", b"00000000000000000000000000000000"),
	(b"01000010001101001011100001010010", b"11000000100001100110011001101000"), -- -49.38 + 45.18 = -4.2
	(b"11000010101110000001010001111011", b"00000000000000000000000000000000"),
	(b"11000010000111011000111101011100", b"11000011000000110110111000010100"), -- -92.04 + -39.39 = -131.43
	(b"01000010011100110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100111000111101011100001", b"01000010001001010010100011110110"), -- 60.85 + -19.56 = 41.29
	(b"11000010100100001101011100001010", b"00000000000000000000000000000000"),
	(b"01000010110000001101000111101100", b"01000001101111111110101110001000"), -- -72.42 + 96.41 = 23.99
	(b"11000001001100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010000001010000000000000000", b"11000010001100010111101011100001"), -- -11.12 + -33.25 = -44.37
	(b"11000001111010000011110101110001", b"00000000000000000000000000000000"),
	(b"11000010000000010011110101110001", b"11000010011101010101110000101010"), -- -29.03 + -32.31 = -61.34
	(b"11000010011101000111000010100100", b"00000000000000000000000000000000"),
	(b"01000010110000100001010001111011", b"01000010000011111011100001010010"), -- -61.11 + 97.04 = 35.93
	(b"01000010001011000001111010111000", b"00000000000000000000000000000000"),
	(b"11000010100000100111010111000011", b"11000001101100011001100110011100"), -- 43.03 + -65.23 = -22.2
	(b"01000010000010000101110000101001", b"00000000000000000000000000000000"),
	(b"11000010000111010011001100110011", b"11000000101001101011100001010000"), -- 34.09 + -39.3 = -5.21
	(b"11000010101110000010111000010100", b"00000000000000000000000000000000"),
	(b"11000000110100010100011110101110", b"11000010110001010100001010001111"), -- -92.09 + -6.54 = -98.63
	(b"11000001111101000001010001111011", b"00000000000000000000000000000000"),
	(b"11000010000011100001111010111000", b"11000010100001000001010001111011"), -- -30.51 + -35.53 = -66.04
	(b"01000010010001000010100011110110", b"00000000000000000000000000000000"),
	(b"11000010011001000101000111101100", b"11000001000000001010001111011000"), -- 49.04 + -57.08 = -8.04
	(b"11000001101000110000101000111101", b"00000000000000000000000000000000"),
	(b"11000001101011000101000111101100", b"11000010001001111010111000010100"), -- -20.38 + -21.54 = -41.92
	(b"01000010100010001101011100001010", b"00000000000000000000000000000000"),
	(b"11000010011110111111010111000011", b"01000000101011011100001010001000"), -- 68.42 + -62.99 = 5.43
	(b"11000000111011000010100011110110", b"00000000000000000000000000000000"),
	(b"11000001101001111100001010001111", b"11000001111000101100110011001100"), -- -7.38 + -20.97 = -28.35
	(b"11000010110000100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000011100011110101110000101", b"11000010101110101010111000010101"), -- -97.12 + 3.78 = -93.34
	(b"11000010000110010001111010111000", b"00000000000000000000000000000000"),
	(b"11000001001111011110101110000101", b"11000010010010001001100110011001"), -- -38.28 + -11.87 = -50.15
	(b"11000001110110101111010111000011", b"00000000000000000000000000000000"),
	(b"11000010101110010101000111101100", b"11000010111100000000111101011101"), -- -27.37 + -92.66 = -120.03
	(b"10111111111000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010101010111011100001010010", b"01000010101010000011001100110011"), -- -1.76 + 85.86 = 84.1
	(b"01000010001100100000101000111101", b"00000000000000000000000000000000"),
	(b"01000001110010111010111000010100", b"01000010100010111111000010100100"), -- 44.51 + 25.46 = 69.97
	(b"11000001010000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000010100010001000101000111101", b"11000010101000001001111010111000"), -- -12.04 + -68.27 = -80.31
	(b"01000010001111010101000111101100", b"00000000000000000000000000000000"),
	(b"11000010101010100010001111010111", b"11000010000101101111010111000010"), -- 47.33 + -85.07 = -37.74
	(b"11000010001110110001010001111011", b"00000000000000000000000000000000"),
	(b"01000001011110000010100011110110", b"11000001111110100001010001111011"), -- -46.77 + 15.51 = -31.26
	(b"01000010101111010011100001010010", b"00000000000000000000000000000000"),
	(b"11000000111100011110101110000101", b"01000010101011100001100110011010"), -- 94.61 + -7.56 = 87.05
	(b"01000000101100000101000111101100", b"00000000000000000000000000000000"),
	(b"11000010010111100011001100110011", b"11000010010010000010100011110110"), -- 5.51 + -55.55 = -50.04
	(b"11000010001101010010100011110110", b"00000000000000000000000000000000"),
	(b"01000001100010100010100011110110", b"11000001111000000010100011110110"), -- -45.29 + 17.27 = -28.02
	(b"11000010100100011101011100001010", b"00000000000000000000000000000000"),
	(b"01000010000000010101110000101001", b"11000010001000100101000111101011"), -- -72.92 + 32.34 = -40.58
	(b"01000001110111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001010011100110011001101", b"01000010100011000100110011001101"), -- 27.7 + 42.45 = 70.15
	(b"11000010100001110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100010100011110101110001", b"11000010101010011111010111000010"), -- -67.7 + -17.28 = -84.98
	(b"11000000001101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000001101111010111000011", b"11000010000100100101110000101001"), -- -2.85 + -33.74 = -36.59
	(b"01000000101010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000010010100010110011001100110", b"01000010011001100111000010100100"), -- 5.26 + 52.35 = 57.61
	(b"01000001111001111110101110000101", b"00000000000000000000000000000000"),
	(b"11000001111010010001111010111000", b"10111110000110011001100110000000"), -- 28.99 + -29.14 = -0.15
	(b"11000001100111111110101110000101", b"00000000000000000000000000000000"),
	(b"01000010101000001101011100001010", b"01000010011100011011100001010010"), -- -19.99 + 80.42 = 60.43
	(b"11000010100011100010001111010111", b"00000000000000000000000000000000"),
	(b"01000010010010101111010111000011", b"11000001101000101010001111010110"), -- -71.07 + 50.74 = -20.33
	(b"11000010011101111110101110000101", b"00000000000000000000000000000000"),
	(b"11000010001100001010111000010100", b"11000010110101000100110011001100"), -- -61.98 + -44.17 = -106.15
	(b"01000010101111000101110000101001", b"00000000000000000000000000000000"),
	(b"01000010010110001000111101011100", b"01000011000101000101000111101100"), -- 94.18 + 54.14 = 148.32
	(b"11000010101011100010001111010111", b"00000000000000000000000000000000"),
	(b"01000010001011001000010100011111", b"11000010001011111100001010001111"), -- -87.07 + 43.13 = -43.94
	(b"01000010011111110111101011100001", b"00000000000000000000000000000000"),
	(b"11000010011100111110101110000101", b"01000000001110001111010111000000"), -- 63.87 + -60.98 = 2.89
	(b"11000010110000000111010111000011", b"00000000000000000000000000000000"),
	(b"11000010001100111000111101011100", b"11000011000011010001111010111000"), -- -96.23 + -44.89 = -141.12
	(b"11000010000001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100111010101110000101001", b"11000010111000000101110000101001"), -- -33.5 + -78.68 = -112.18
	(b"11000010010000011010001111010111", b"00000000000000000000000000000000"),
	(b"11000000100011000111101011100001", b"11000010010100110011001100110011"), -- -48.41 + -4.39 = -52.8
	(b"01000010001000011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010110000010111010111000011", b"11000010011000010000000000000001"), -- 40.48 + -96.73 = -56.25
	(b"01000000010001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000010101101001000010100011111", b"01000010101110101100001010010000"), -- 3.12 + 90.26 = 93.38
	(b"11000001101010100010100011110110", b"00000000000000000000000000000000"),
	(b"11000010110001101011100001010010", b"11000010111100010100001010010000"), -- -21.27 + -99.36 = -120.63
	(b"01000001100001101010001111010111", b"00000000000000000000000000000000"),
	(b"11000010101100010110000101001000", b"11000010100011111011100001010010"), -- 16.83 + -88.69 = -71.86
	(b"01000010000101101110101110000101", b"00000000000000000000000000000000"),
	(b"01000010000001110110011001100110", b"01000010100011110010100011110110"), -- 37.73 + 33.85 = 71.58
	(b"01000010100001010101011100001010", b"00000000000000000000000000000000"),
	(b"11000010101111010000000000000000", b"11000001110111101010001111011000"), -- 66.67 + -94.5 = -27.83
	(b"01000010001010100100011110101110", b"00000000000000000000000000000000"),
	(b"01000010101000111100011110101110", b"01000010111110001110101110000101"), -- 42.57 + 81.89 = 124.46
	(b"11000010011011000010100011110110", b"00000000000000000000000000000000"),
	(b"11000010000011000001010001111011", b"11000010101111000001111010111000"), -- -59.04 + -35.02 = -94.06
	(b"11000001100100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001011010100011110101110001", b"11000010000001000101110000101001"), -- -18.45 + -14.64 = -33.09
	(b"01000010101001000000101000111101", b"00000000000000000000000000000000"),
	(b"11000010100000011000000000000000", b"01000001100010100010100011110100"), -- 82.02 + -64.75 = 17.27
	(b"11000010101010001011100001010010", b"00000000000000000000000000000000"),
	(b"11000010001110110010100011110110", b"11000011000000110010011001100110"), -- -84.36 + -46.79 = -131.15
	(b"11000010100111011000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001101010101000111101100", b"11000010111110000010100011110110"), -- -78.75 + -45.33 = -124.08
	(b"01000010100010111000101000111101", b"00000000000000000000000000000000"),
	(b"01000000100100001111010111000011", b"01000010100101001001100110011001"), -- 69.77 + 4.53 = 74.3
	(b"01000010100100000001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001010010010100011110110", b"01000010111001001010111000010101"), -- 72.05 + 42.29 = 114.34
	(b"01000010100010100101011100001010", b"00000000000000000000000000000000"),
	(b"11000001111111100110011001100110", b"01000010000101010111101011100001"), -- 69.17 + -31.8 = 37.37
	(b"01000010101001000100011110101110", b"00000000000000000000000000000000"),
	(b"11000010010011010010100011110110", b"01000001111101101100110011001100"), -- 82.14 + -51.29 = 30.85
	(b"01000001111111100010100011110110", b"00000000000000000000000000000000"),
	(b"11000010001011011110101110000101", b"11000001001110110101110000101000"), -- 31.77 + -43.48 = -11.71
	(b"01000010110000100101110000101001", b"00000000000000000000000000000000"),
	(b"11000010001000010000000000000000", b"01000010011000111011100001010010"), -- 97.18 + -40.25 = 56.93
	(b"01000010100010100110000101001000", b"00000000000000000000000000000000"),
	(b"11000010000100110011110101110001", b"01000010000000011000010100011111"), -- 69.19 + -36.81 = 32.38
	(b"11000010010010001011100001010010", b"00000000000000000000000000000000"),
	(b"11000010100011010111000010100100", b"11000010111100011100110011001101"), -- -50.18 + -70.72 = -120.9
	(b"11000001110001100011110101110001", b"00000000000000000000000000000000"),
	(b"11000001010000001100110011001101", b"11000010000100110101000111101100"), -- -24.78 + -12.05 = -36.83
	(b"01000010101111010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000111010110011001100110", b"01000010010111001001100110011010"), -- 94.5 + -39.35 = 55.15
	(b"01000010000011101110101110000101", b"00000000000000000000000000000000"),
	(b"01000010100001000000101000111101", b"01000010110010111000000000000000"), -- 35.73 + 66.02 = 101.75
	(b"11000010101011011101011100001010", b"00000000000000000000000000000000"),
	(b"11000010101001010111010111000011", b"11000011001010011010011001100110"), -- -86.92 + -82.73 = -169.65
	(b"11000010100101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111101101011100001010", b"11000001100100100101000111101100"), -- -74 + 55.71 = -18.29
	(b"11000010100101100111101011100001", b"00000000000000000000000000000000"),
	(b"11000000100101011100001010001111", b"11000010100111111101011100001010"), -- -75.24 + -4.68 = -79.92
	(b"01000000100110111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010101011000011110101110001", b"01000010101101011111101011100010"), -- 4.87 + 86.12 = 90.99
	(b"01000010011011001010001111010111", b"00000000000000000000000000000000"),
	(b"01000010100010011100110011001101", b"01000011000000000000111101011100"), -- 59.16 + 68.9 = 128.06
	(b"01000010001100100100011110101110", b"00000000000000000000000000000000"),
	(b"01000010001001000100011110101110", b"01000010101010110100011110101110"), -- 44.57 + 41.07 = 85.64
	(b"11000010001001111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101100100010001111010111", b"11000011000000110000010100011111"), -- -41.95 + -89.07 = -131.02
	(b"01000010100100111000111101011100", b"00000000000000000000000000000000"),
	(b"11000010000000110001010001111011", b"01000010001001000000101000111101"), -- 73.78 + -32.77 = 41.01
	(b"01000010000000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011101100011001100110011", b"11000001111001010011001100110010"), -- 32.9 + -61.55 = -28.65
	(b"10111111100000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010001110111111010111000011", b"01000010001101111110101110000110"), -- -1.01 + 46.99 = 45.98
	(b"01000010101110101001111010111000", b"00000000000000000000000000000000"),
	(b"11000010000101010001010001111011", b"01000010011000000010100011110101"), -- 93.31 + -37.27 = 56.04
	(b"11000010010001111011100001010010", b"00000000000000000000000000000000"),
	(b"01000001101100011100001010001111", b"11000001110111011010111000010101"), -- -49.93 + 22.22 = -27.71
	(b"11000010110000110111101011100001", b"00000000000000000000000000000000"),
	(b"11000010101010011111000010100100", b"11000011001101101011010111000010"), -- -97.74 + -84.97 = -182.71
	(b"01000001011011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111110111101011100001010", b"11000001100001001010001111010111"), -- 14.9 + -31.48 = -16.58
	(b"11000010000101001111010111000011", b"00000000000000000000000000000000"),
	(b"01000001011110101011100001010010", b"11000001101011001000111101011101"), -- -37.24 + 15.67 = -21.57
	(b"01000010100000111001010001111011", b"00000000000000000000000000000000"),
	(b"10111110011010111000010100011111", b"01000010100000110001111010111000"), -- 65.79 + -0.23 = 65.56
	(b"01000010110001110110101110000101", b"00000000000000000000000000000000"),
	(b"01000001000100010001111010111000", b"01000010110110011000111101011100"), -- 99.71 + 9.07 = 108.78
	(b"11000010100110010010001111010111", b"00000000000000000000000000000000"),
	(b"01000001110111011000010100011111", b"11000010010000111000010100011110"), -- -76.57 + 27.69 = -48.88
	(b"11000010100101111011100001010010", b"00000000000000000000000000000000"),
	(b"11000001100110000000000000000000", b"11000010101111011011100001010010"), -- -75.86 + -19 = -94.86
	(b"11000010100111000011100001010010", b"00000000000000000000000000000000"),
	(b"11000010100011110001010001111011", b"11000011000101011010011001100110"), -- -78.11 + -71.54 = -149.65
	(b"01000001010011000101000111101100", b"00000000000000000000000000000000"),
	(b"01000001011000110101110000101001", b"01000001110101111101011100001010"), -- 12.77 + 14.21 = 26.98
	(b"01000010100101001011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000000101110101110000101", b"01000010110101100010100011110110"), -- 74.35 + 32.73 = 107.08
	(b"11000010101011011100011110101110", b"00000000000000000000000000000000"),
	(b"01000001100100101010001111010111", b"11000010100010010001111010111000"), -- -86.89 + 18.33 = -68.56
	(b"11000010000011110000101000111101", b"00000000000000000000000000000000"),
	(b"01000001000101110000101000111101", b"11000001110100101000111101011100"), -- -35.76 + 9.44 = -26.32
	(b"11000001111111010001111010111000", b"00000000000000000000000000000000"),
	(b"11000010101111011100011110101110", b"11000010111111010000111101011100"), -- -31.64 + -94.89 = -126.53
	(b"11000010101111101101110000101001", b"00000000000000000000000000000000"),
	(b"01000010101101011101000111101100", b"11000000100100001010001111010000"), -- -95.43 + 90.91 = -4.52
	(b"11000001110000111010111000010100", b"00000000000000000000000000000000"),
	(b"01000010010111100001111010111000", b"01000001111110001000111101011100"), -- -24.46 + 55.53 = 31.07
	(b"11000010011000001110000101001000", b"00000000000000000000000000000000"),
	(b"11000010100010010000000000000000", b"11000010111110010111000010100100"), -- -56.22 + -68.5 = -124.72
	(b"01000010101100101000010100011111", b"00000000000000000000000000000000"),
	(b"11000010110000001111000010100100", b"11000000111001101011100001010000"), -- 89.26 + -96.47 = -7.21
	(b"11000010011100010000101000111101", b"00000000000000000000000000000000"),
	(b"01000010010111011100110011001101", b"11000000100110011110101110000000"), -- -60.26 + 55.45 = -4.81
	(b"01000001101011101111010111000011", b"00000000000000000000000000000000"),
	(b"01000010000011000100011110101110", b"01000010011000111100001010010000"), -- 21.87 + 35.07 = 56.94
	(b"01000010100010100010111000010100", b"00000000000000000000000000000000"),
	(b"01000010101001100110101110000101", b"01000011000110000100110011001100"), -- 69.09 + 83.21 = 152.3
	(b"11000001111111111100001010001111", b"00000000000000000000000000000000"),
	(b"01000010101100001111010111000011", b"01000010011000100000101000111110"), -- -31.97 + 88.48 = 56.51
	(b"01000010010111011110101110000101", b"00000000000000000000000000000000"),
	(b"01000010100001111101011100001010", b"01000010111101101100110011001100"), -- 55.48 + 67.92 = 123.4
	(b"11000010010000110001010001111011", b"00000000000000000000000000000000"),
	(b"01000010001010111010111000010100", b"11000000101110110011001100111000"), -- -48.77 + 42.92 = -5.85
	(b"11000010011010101000111101011100", b"00000000000000000000000000000000"),
	(b"11000010000110110111101011100001", b"11000010110000110000010100011110"), -- -58.64 + -38.87 = -97.51
	(b"11000010010011011000111101011100", b"00000000000000000000000000000000"),
	(b"01000010011111110011110101110001", b"01000001010001101011100001010100"), -- -51.39 + 63.81 = 12.42
	(b"01000010100100110011100001010010", b"00000000000000000000000000000000"),
	(b"01000001011101001010001111010111", b"01000010101100011100110011001101"), -- 73.61 + 15.29 = 88.9
	(b"01000010011011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110110110001111010111000", b"01000010000000000000101000111110"), -- 59.4 + -27.39 = 32.01
	(b"11000010000001101101011100001010", b"00000000000000000000000000000000"),
	(b"01000001111010111000010100011111", b"11000000100010001010001111010100"), -- -33.71 + 29.44 = -4.27
	(b"11000010100111011011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001100101110000101001000", b"11000010000010001000010100011110"), -- -78.85 + 44.72 = -34.13
	(b"01000001100010101000111101011100", b"00000000000000000000000000000000"),
	(b"01000001101110011001100110011010", b"01000010001000100001010001111011"), -- 17.32 + 23.2 = 40.52
	(b"11000010001011001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010110110001010001111011", b"01000001001110011110101110000100"), -- -43.15 + 54.77 = 11.62
	(b"11000010001000100111101011100001", b"00000000000000000000000000000000"),
	(b"01000001111000000111101011100001", b"11000001010010001111010111000010"), -- -40.62 + 28.06 = -12.56
	(b"11000010110000010101000111101100", b"00000000000000000000000000000000"),
	(b"11000010100001001000010100011111", b"11000011001000101110101110000110"), -- -96.66 + -66.26 = -162.92
	(b"01000010100001010010001111010111", b"00000000000000000000000000000000"),
	(b"01000010000011111000111101011100", b"01000010110011001110101110000101"), -- 66.57 + 35.89 = 102.46
	(b"11000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000010100111110100110011001101", b"01000010100101110101011100001010"), -- -3.98 + 79.65 = 75.67
	(b"11000010101011000100001010001111", b"00000000000000000000000000000000"),
	(b"01000010001101010110011001100110", b"11000010001000110001111010111000"), -- -86.13 + 45.35 = -40.78
	(b"11000010100110100001010001111011", b"00000000000000000000000000000000"),
	(b"01000010101100110011001100110011", b"01000001010010001111010111000000"), -- -77.04 + 89.6 = 12.56
	(b"11000001111110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001101010111001100110011010", b"11000010010100110011110101110001"), -- -31.36 + -21.45 = -52.81
	(b"11000010110001010100001010001111", b"00000000000000000000000000000000"),
	(b"11000001110110001000111101011100", b"11000010111110110110011001100110"), -- -98.63 + -27.07 = -125.7
	(b"11000010100111010111010111000011", b"00000000000000000000000000000000"),
	(b"11000001100000111100001010001111", b"11000010101111100110011001100111"), -- -78.73 + -16.47 = -95.2
	(b"11000001110100111100001010001111", b"00000000000000000000000000000000"),
	(b"11000010100000000101011100001010", b"11000010101101010100011110101110"), -- -26.47 + -64.17 = -90.64
	(b"11000010010011011110101110000101", b"00000000000000000000000000000000"),
	(b"11000010110001001011001100110011", b"11000011000101011101010001111011"), -- -51.48 + -98.35 = -149.83
	(b"11000010000001011010001111010111", b"00000000000000000000000000000000"),
	(b"11000010000100011010111000010100", b"11000010100010111010100011110110"), -- -33.41 + -36.42 = -69.83
	(b"11000010000110100100011110101110", b"00000000000000000000000000000000"),
	(b"11000001100110011010111000010100", b"11000010011001110001111010111000"), -- -38.57 + -19.21 = -57.78
	(b"11000001111111111110101110000101", b"00000000000000000000000000000000"),
	(b"01000001110011011100001010001111", b"11000000110010001010001111011000"), -- -31.99 + 25.72 = -6.27
	(b"11000010101011010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100000101110000101001000", b"11000010110011011011100001010010"), -- -86.5 + -16.36 = -102.86
	(b"11000010010111101000111101011100", b"00000000000000000000000000000000"),
	(b"11000010011111001111010111000011", b"11000010111011011100001010010000"), -- -55.64 + -63.24 = -118.88
	(b"11000010000011110001111010111000", b"00000000000000000000000000000000"),
	(b"01000010011100000111101011100001", b"01000001110000101011100001010010"), -- -35.78 + 60.12 = 24.34
	(b"01000010010010010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111100001010001111011", b"01000010110100111000101000111110"), -- 50.25 + 55.52 = 105.77
	(b"11000010011010011000111101011100", b"00000000000000000000000000000000"),
	(b"11000001011010001111010111000011", b"11000010100100011110011001100110"), -- -58.39 + -14.56 = -72.95
	(b"01000010011100100111000010100100", b"00000000000000000000000000000000"),
	(b"01000010001101110110011001100110", b"01000010110101001110101110000101"), -- 60.61 + 45.85 = 106.46
	(b"11000010000000111110000101001000", b"00000000000000000000000000000000"),
	(b"11000010101100100111000010100100", b"11000010111101000110000101001000"), -- -32.97 + -89.22 = -122.19
	(b"11000001100110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010110000000110101110000101", b"11000010111001101011100001010010"), -- -19.15 + -96.21 = -115.36
	(b"11000010101110111101110000101001", b"00000000000000000000000000000000"),
	(b"01000010001110111100110011001101", b"11000010001110111110101110000101"), -- -93.93 + 46.95 = -46.98
	(b"11000010011010111011100001010010", b"00000000000000000000000000000000"),
	(b"11000010101011000010001111010111", b"11000011000100010000000000000000"), -- -58.93 + -86.07 = -145
	(b"01000001101011111110101110000101", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000001111000111110101110000101"), -- 21.99 + 6.5 = 28.49
	(b"01000000111000001111010111000011", b"00000000000000000000000000000000"),
	(b"11000001011101000101000111101100", b"11000001000000111101011100001010"), -- 7.03 + -15.27 = -8.24
	(b"11000010100111101100011110101110", b"00000000000000000000000000000000"),
	(b"01000001101000111110101110000101", b"11000010011010111001100110011010"), -- -79.39 + 20.49 = -58.9
	(b"01000010000010010010100011110110", b"00000000000000000000000000000000"),
	(b"11000010101110000111010111000011", b"11000010011001111100001010010000"), -- 34.29 + -92.23 = -57.94
	(b"11000001001011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000010100000111000111101011100", b"01000010010110111001100110011001"), -- -10.88 + 65.78 = 54.9
	(b"11000010100000001010100011110110", b"00000000000000000000000000000000"),
	(b"01000010101010011110000101001000", b"01000001101001001110000101001000"), -- -64.33 + 84.94 = 20.61
	(b"11000010010101110100011110101110", b"00000000000000000000000000000000"),
	(b"11000010100000101101000111101100", b"11000010111011100111010111000011"), -- -53.82 + -65.41 = -119.23
	(b"01000000100010010100011110101110", b"00000000000000000000000000000000"),
	(b"01000010001011111010111000010100", b"01000010010000001101011100001010"), -- 4.29 + 43.92 = 48.21
	(b"11000010101011010010001111010111", b"00000000000000000000000000000000"),
	(b"11000010101100101001100110011010", b"11000011001011111101111010111000"), -- -86.57 + -89.3 = -175.87
	(b"01000010000110101010111000010100", b"00000000000000000000000000000000"),
	(b"01000010011110011001100110011010", b"01000010110010100010001111010111"), -- 38.67 + 62.4 = 101.07
	(b"11000001010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110111110101110000101001000", b"11000001010101110011001100110011"), -- -12.96 + -0.49 = -13.45
	(b"01000010100100100110101110000101", b"00000000000000000000000000000000"),
	(b"11000010100000010010100011110110", b"01000001000010100001010001111000"), -- 73.21 + -64.58 = 8.63
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000011111010111000010100", b"01000000101101011100001010001110"), -- -3.3 + 8.98 = 5.68
	(b"11000010010000010001111010111000", b"00000000000000000000000000000000"),
	(b"11000010110001010101000111101100", b"11000011000100101111000010100100"), -- -48.28 + -98.66 = -146.94
	(b"01000001101101101010001111010111", b"00000000000000000000000000000000"),
	(b"01000010010100000101000111101100", b"01000010100101011101000111101100"), -- 22.83 + 52.08 = 74.91
	(b"01000001101000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000001101011111101011100001010", b"10111111110101000111101011100000"), -- 20.32 + -21.98 = -1.66
	(b"11000000111001101011100001010010", b"00000000000000000000000000000000"),
	(b"01000010100011000111010111000011", b"01000010011111000001010001111100"), -- -7.21 + 70.23 = 63.02
	(b"11000010101100111011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011101000111101011100", b"11000010110001011000010100011110"), -- -89.85 + -8.91 = -98.76
	(b"01000001011100100011110101110001", b"00000000000000000000000000000000"),
	(b"11000001110010000101000111101100", b"11000001000111100110011001100111"), -- 15.14 + -25.04 = -9.9
	(b"01000010000111001001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000001010001111010111000", b"01000010000110101000010100011111"), -- 39.15 + -0.52 = 38.63
	(b"01000010011011111011100001010010", b"00000000000000000000000000000000"),
	(b"01000010101010001110011001100110", b"01000011000100000110000101001000"), -- 59.93 + 84.45 = 144.38
	(b"01000010100100001111010111000011", b"00000000000000000000000000000000"),
	(b"01000001000101000010100011110110", b"01000010101000110111101011100010"), -- 72.48 + 9.26 = 81.74
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000100010101110000101001000", b"01000000011011101011100001010010"), -- -0.61 + 4.34 = 3.73
	(b"11000010101011101011110101110001", b"00000000000000000000000000000000"),
	(b"01000010110000110001010001111011", b"01000001001000101011100001010000"), -- -87.37 + 97.54 = 10.17
	(b"11000001101001100111101011100001", b"00000000000000000000000000000000"),
	(b"01000010100111011010001111010111", b"01000010011010000000101000111110"), -- -20.81 + 78.82 = 58.01
	(b"11000001101100000111101011100001", b"00000000000000000000000000000000"),
	(b"11000010100000000000000000000000", b"11000010101011000001111010111000"), -- -22.06 + -64 = -86.06
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010000001001100110011010", b"11000010011000110110011001100111"), -- -8.7 + -48.15 = -56.85
	(b"11000001000001111101011100001010", b"00000000000000000000000000000000"),
	(b"01000010100111010101110000101001", b"01000010100011000110000101001000"), -- -8.49 + 78.68 = 70.19

	(b"01000000100001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101010101110000101001000", b"10111111100110000101000111101100"), -- 4.15 + -5.34 = -1.19
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000011110101110000101", b"11000000110001000010100011110110"), -- -2.6 + -3.53 = -6.13
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"00111111001100001010001111010111"), -- 0.22 + 0.47 = 0.69
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000001000111000000000000000000", b"11000001000111001111010111000011"), -- -0.06 + -9.75 = -9.81
	(b"01000000110011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000101111110000101000111101", b"01000001010001101000111101011100"), -- 6.44 + 5.97 = 12.41
	(b"01000001000110101011100001010010", b"00000000000000000000000000000000"),
	(b"11000001000010110000101000111101", b"00111111011110101110000101010000"), -- 9.67 + -8.69 = 0.98
	(b"11000000111001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000011000111101011100001010", b"11000001001011001100110011001100"), -- -7.24 + -3.56 = -10.8
	(b"01000001000001010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111110111010111000010100100", b"01000001001000001111010111000010"), -- 8.33 + 1.73 = 10.06
	(b"11000000110011111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110100000000000000000000000", b"11000000110101111010111000010100"), -- -6.49 + -0.25 = -6.74
	(b"01000001000000110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000111000101110000101001000", b"00111111100011001100110011001000"), -- 8.19 + -7.09 = 1.1
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000001000001000101000111101100", b"11000000111111010001111010111001"), -- 0.36 + -8.27 = -7.91
	(b"01000000000001000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000010010000101000111101100", b"10111111100001111010111000010110"), -- 2.07 + -3.13 = -1.06
	(b"00111111100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111110111101011100001010", b"11000000110101110000101000111101"), -- 1.15 + -7.87 = -6.72
	(b"01000000100000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000110110001111010111000011", b"11000000001011001100110011001110"), -- 4.08 + -6.78 = -2.7
	(b"00111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000110100011001100110011010", b"01000000111011000111101011100010"), -- 0.84 + 6.55 = 7.39
	(b"10111111100001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"10111111000100011110101110000100"), -- -1.04 + 0.47 = -0.57
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111001110101110000101001", b"11000001001000111010111000010100"), -- -3 + -7.23 = -10.23
	(b"11000001000110101000111101011100", b"00000000000000000000000000000000"),
	(b"01000001000000110000101000111101", b"10111111101111000010100011111000"), -- -9.66 + 8.19 = -1.47
	(b"11000001000001000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000110111000010100011110101"), -- -8.28 + 1.4 = -6.88
	(b"01000001000011111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"01000000101111000111101011100001"), -- 8.99 + -3.1 = 5.89
	(b"01000000001011000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000101101000010100011110110", b"01000001000001010001111010111000"), -- 2.69 + 5.63 = 8.32
	(b"10111111100100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000001000010100001010001111011", b"11000001000111000010100011110110"), -- -1.13 + -8.63 = -9.76
	(b"10111111100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100110001010001111010111", b"11000000101110100011110101110000"), -- -1.05 + -4.77 = -5.82
	(b"11000000100000100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000000110101110000101001000", b"11000000110011111010111000010101"), -- -4.07 + -2.42 = -6.49
	(b"01000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000111010010100011110101110", b"01000001001001000010100011110110"), -- 2.97 + 7.29 = 10.26
	(b"11000000000100010100011110101110", b"00000000000000000000000000000000"),
	(b"01000001000000100011110101110001", b"01000000101110111101011100001011"), -- -2.27 + 8.14 = 5.87
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000100100011110101110001", b"01000001000101110000101000111110"), -- 0.3 + 9.14 = 9.44
	(b"01000000010000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000001000101000010100011110110", b"01000001010001001100110011001101"), -- 3.04 + 9.26 = 12.3
	(b"01000000110011000010100011110110", b"00000000000000000000000000000000"),
	(b"11000001000010101000111101011100", b"11000000000100011110101110000100"), -- 6.38 + -8.66 = -2.28
	(b"11000000110010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010101111010111000010100", b"11000000001111001100110011001110"), -- -6.32 + 3.37 = -2.95
	(b"00111111101010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000001000100110101110000101001", b"11000000111111000010100011110110"), -- 1.33 + -9.21 = -7.88
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000101000010100011110101110", b"01000000101101101011100001010010"), -- 0.67 + 5.04 = 5.71
	(b"01000000010100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000010010100011110101110001", b"01000000110011010111000010100100"), -- 3.26 + 3.16 = 6.42
	(b"00111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000001000010100110011001100110", b"01000001000011001111010111000010"), -- 0.16 + 8.65 = 8.81
	(b"01000000110110101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000101101110101110000101001"), -- 6.83 + -1.1 = 5.73
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000001000101000111101100", b"11000000101110001010001111011000"), -- 2.5 + -8.27 = -5.77
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"00111111000111000010100011110110"), -- 0.54 + 0.07 = 0.61
	(b"11000000000000001010001111010111", b"00000000000000000000000000000000"),
	(b"01000001000111011100001010001111", b"01000000111110110011001100110010"), -- -2.01 + 9.86 = 7.85
	(b"00111111101011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000100110000101000111101100", b"01000000110001000010100011110110"), -- 1.37 + 4.76 = 6.13
	(b"01000000111111110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"01000001000001011001100110011001"), -- 7.97 + 0.38 = 8.35
	(b"01000001000101010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"01000000100001110000101000111101"), -- 9.32 + -5.1 = 4.22
	(b"01000000101101010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"01000000101110110011001100110011"), -- 5.66 + 0.19 = 5.85
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101111000010100011111", b"01000001010111011110101110000110"), -- 4.4 + 9.47 = 13.87
	(b"01000000110111110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"01000000101111111010111000010100"), -- 6.98 + -0.99 = 5.99
	(b"11000000000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000100100110011001100110", b"11000001001100110011001100110011"), -- -2.05 + -9.15 = -11.2
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000000011100001010001111011", b"11000000000111010111000010100100"), -- -0.24 + -2.22 = -2.46
	(b"11000000010000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011011100001010001111011", b"11000000011111110101110000101001"), -- -3.06 + -0.93 = -3.99
	(b"11000000101011000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000000011100001010001111011", b"11000000111100110011001100110100"), -- -5.38 + -2.22 = -7.6
	(b"01000001000011011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111110101011100001010001111", b"01000001001010001010001111010111"), -- 8.87 + 1.67 = 10.54
	(b"01000001000101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110011000111101011100001", b"01000001011110111101011100001010"), -- 9.35 + 6.39 = 15.74
	(b"01000000100000001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000111010101000111101011100", b"01000001001101011100001010010000"), -- 4.03 + 7.33 = 11.36
	(b"10111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111111010111000010100100", b"11000000001000011110101110000101"), -- -0.55 + -1.98 = -2.53
	(b"11000000111111011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000100001101011100001010010", b"11000001010000100011110101110000"), -- -7.93 + -4.21 = -12.14
	(b"11000001000010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000001000101111000010100011111", b"00111111010101000111101011100000"), -- -8.64 + 9.47 = 0.83
	(b"10111111101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000011001011100001010001111", b"11000000100110111101011100001010"), -- -1.28 + -3.59 = -4.87
	(b"01000000100001010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000001000111000101000111101100"), -- 4.17 + 5.6 = 9.77
	(b"11000000100000101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000010111000010100011110110", b"10111111001001100110011001101000"), -- -4.09 + 3.44 = -0.65
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001000011010111000010100100"), -- 0.86 + -9.7 = -8.84
	(b"11000000010101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100010111101011100001010", b"11000000111101110000101000111101"), -- -3.35 + -4.37 = -7.72
	(b"01000000101111000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000011000011110101110000101", b"01000001000101101011100001010010"), -- 5.89 + 3.53 = 9.42
	(b"11000000111001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000100001010111000010100100", b"11000001001101100011110101110000"), -- -7.22 + -4.17 = -11.39
	(b"00111111100110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000001010111000010100011111", b"01000000011110001111010111000011"), -- 1.21 + 2.68 = 3.89
	(b"01000000000000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000110110001010001111010111", b"01000001000011010100011110101110"), -- 2.06 + 6.77 = 8.83
	(b"11000001000110001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000101100111000010100011111", b"11000000011111001100110011001110"), -- -9.56 + 5.61 = -3.95
	(b"11000001000000110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000111110100011110101110001", b"11000001100000000011110101110001"), -- -8.21 + -7.82 = -16.03
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110001110101110000101001", b"01000001001011101110000101001000"), -- 4.7 + 6.23 = 10.93
	(b"10111111111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110111000010100011111", b"00111111001011100001010001111100"), -- -1.75 + 2.43 = 0.68
	(b"01000001000001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000101111101011100001010", b"10111111100100011110101110000000"), -- 8.35 + -9.49 = -1.14
	(b"01000000110111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000110110110011001100110011", b"00111100111101011100001100000000"), -- 6.88 + -6.85 = 0.0300002
	(b"10111111111111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000000100001110000101000111101"), -- -1.98 + 6.2 = 4.22
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111111011100001010001111011", b"00111111101010001111010111000010"), -- -0.54 + 1.86 = 1.32
	(b"11000000110010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000101001011100001010001111", b"10111111100100011110101110001000"), -- -6.32 + 5.18 = -1.14
	(b"11000000111011010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"11000001000001010100011110101110"), -- -7.42 + -0.91 = -8.33
	(b"11000000110001101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000110101000010100011110110", b"11000001010011010111000010100100"), -- -6.21 + -6.63 = -12.84
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111010101000111101011100010"), -- 0.37 + -1.2 = -0.83
	(b"01000000000000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"00111111111010100011110101110000"), -- 2.05 + -0.22 = 1.83
	(b"11000001000001011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000000100011110101110000101", b"11000001001010100011110101110000"), -- -8.36 + -2.28 = -10.64
	(b"01000000110111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000100101100001010001111011", b"01000001001110010001111010111000"), -- 6.88 + 4.69 = 11.57
	(b"10111111111001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000001000110011100001010001111", b"11000001001101100110011001100110"), -- -1.79 + -9.61 = -11.4
	(b"11000000101101101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000100110000000000000000000", b"10111111011101011100001010010000"), -- -5.71 + 4.75 = -0.96
	(b"11000000111011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111000100011110101110000101", b"11000000110110111101011100001010"), -- -7.44 + 0.57 = -6.87
	(b"11000000111111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000000111001100110011001101", b"11000001001001011110101110000101"), -- -7.92 + -2.45 = -10.37
	(b"11000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111101111000010100011110101110", b"11000000011101111010111000010101"), -- -3.98 + 0.11 = -3.87
	(b"01000000111110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000011111101011100001010010", b"01000000011100011110101110000110"), -- 7.76 + -3.98 = 3.78
	(b"01000000110101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000001000101100001010001111011", b"01000001100000001100110011001101"), -- 6.72 + 9.38 = 16.1
	(b"10111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000000000110011001100110011", b"00111111101010001111010111000010"), -- -0.73 + 2.05 = 1.32
	(b"00111111101010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"00111111000001010001111010111001"), -- 1.34 + -0.82 = 0.52
	(b"11000001000001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000110111100001010001111011", b"11000001011101000010100011110110"), -- -8.32 + -6.94 = -15.26
	(b"11000000000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100010110011001100110011", b"11000000110110011001100110011010"), -- -2.45 + -4.35 = -6.8
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000001000000000000000000", b"11000001001000001100110011001101"), -- -1.8 + -8.25 = -10.05
	(b"01000000110001000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"10111111000100011110101110000000"), -- 6.13 + -6.7 = -0.57
	(b"11000001000011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111011110101110000101001", b"10111111101111000010100011110100"), -- -8.95 + 7.48 = -1.47
	(b"11000001000110101011100001010010", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001100101010101110000101001"), -- -9.67 + -9 = -18.67
	(b"11000000110100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010101010001111010111000", b"11000001000111011001100110011010"), -- -6.52 + -3.33 = -9.85
	(b"11000000010101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"11000000000110000101000111101011"), -- -3.32 + 0.94 = -2.38
	(b"11000001000100010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000110000111101011100001010", b"11000001011100110101110000101001"), -- -9.09 + -6.12 = -15.21
	(b"01000001000100101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000001001111010111000010100", b"01000000110100010100011110101110"), -- 9.16 + -2.62 = 6.54
	(b"01000000101000100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000110001001100110011001101", b"10111111100010100011110101110000"), -- 5.07 + -6.15 = -1.08
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000001000010100011110110", b"11000001000010000010100011110110"), -- -0.25 + -8.26 = -8.51
	(b"00111111111000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000110000011001100110011010", b"01000000111110101000111101011100"), -- 1.78 + 6.05 = 7.83
	(b"01000000100000101110000101001000", b"00000000000000000000000000000000"),
	(b"01000001000010000101000111101100", b"01000001010010011100001010010000"), -- 4.09 + 8.52 = 12.61
	(b"01000000101011000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000111101010111000010100100", b"01000001010100001111010111000010"), -- 5.39 + 7.67 = 13.06
	(b"11000000001101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000101101010111000010100100", b"01000000001101010001111010111001"), -- -2.84 + 5.67 = 2.83
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000101000111101011100001", b"01000001010101000111101011100001"), -- 4 + 9.28 = 13.28
	(b"11000000011001000111101011100001", b"00000000000000000000000000000000"),
	(b"11000001000001110101110000101001", b"11000001010000000111101011100001"), -- -3.57 + -8.46 = -12.03
	(b"11000000000010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000101101110000101000111101", b"01000000011000110011001100110010"), -- -2.17 + 5.72 = 3.55
	(b"01000000111100111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000101010010100011110101110", b"01000000000101000111101011100010"), -- 7.61 + -5.29 = 2.32
	(b"11000001000000001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000001100010100011110101110", b"11000000101010001010001111010111"), -- -8.04 + 2.77 = -5.27
	(b"11000000011000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000000110001111010111000010101"), -- -3.56 + 9.8 = 6.24
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000001000100001100110011001101", b"11000001001000000010100011110110"), -- -0.96 + -9.05 = -10.01
	(b"01000000101110100011110101110001", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000000001111101011100001010010"), -- 5.82 + -8.8 = -2.98
	(b"01000000101111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111100110101110000101001000", b"01000000100110000000000000000000"), -- 5.96 + -1.21 = 4.75
	(b"11000000110010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000001000000101011100001010010", b"11000001011001110011001100110100"), -- -6.28 + -8.17 = -14.45
	(b"01000000100100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000011000001010001111010111", b"01000001000000000111101011100001"), -- 4.52 + 3.51 = 8.03
	(b"01000000111100111000010100011111", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000001011111001111010111000010"), -- 7.61 + 8.2 = 15.81
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000001000010100001010001111011", b"01000000111110000101000111101100"), -- -0.87 + 8.63 = 7.76
	(b"11000000101001010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000101010000101000111101100", b"11000001001001101110000101001000"), -- -5.17 + -5.26 = -10.43
	(b"11000000100001000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000001111000010100011110110", b"11000000111000100011110101110001"), -- -4.13 + -2.94 = -7.07
	(b"11000000100111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000100101100001010001111011", b"10111110010000101000111101100000"), -- -4.88 + 4.69 = -0.19
	(b"01000000110111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111011100110011001100110011", b"01000000111110111101011100001010"), -- 6.92 + 0.95 = 7.87
	(b"01000000011011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000010011101011100001010010", b"00111111000000101000111101011100"), -- 3.74 + -3.23 = 0.51
	(b"01000000001010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000010111000010100100", b"11000000101011100001010001111011"), -- 2.65 + -8.09 = -5.44
	(b"01000000101011000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000011011100001010001111011", b"01000001000100011100001010001111"), -- 5.39 + 3.72 = 9.11
	(b"11000000000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111100010111000010100011111", b"10111111100100110011001100110011"), -- -2.24 + 1.09 = -1.15
	(b"01000001000001111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"01000001000011000111101011100001"), -- 8.49 + 0.29 = 8.78
	(b"11000001000000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101000111101011100001", b"10111111101101000111101011100100"), -- -8.05 + 6.64 = -1.41
	(b"01000000100110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000101101000111101011100001", b"10111111011000010100011110101000"), -- 4.76 + -5.64 = -0.88
	(b"11000000111000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000110001110000101000111101", b"11000001010101010111000010100100"), -- -7.12 + -6.22 = -13.34
	(b"11000001000010100001010001111011", b"00000000000000000000000000000000"),
	(b"01000001000111011110101110000101", b"00111111100111101011100001010000"), -- -8.63 + 9.87 = 1.24
	(b"11000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000001000000001111010111000011", b"01000000101010000000000000000001"), -- -2.81 + 8.06 = 5.25
	(b"01000000000000011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000101000100011110101110001", b"01000000111000110011001100110100"), -- 2.03 + 5.07 = 7.1
	(b"00111111100001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000110001101011100001010010", b"01000000111010001010001111010111"), -- 1.06 + 6.21 = 7.27
	(b"01000001000101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110000001111010111000011", b"01000000010101000111101011100010"), -- 9.35 + -6.03 = 3.32
	(b"11000000010111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"00111111001101011100001010001100"), -- -3.49 + 4.2 = 0.71
	(b"11000000111000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101000000101000111101100", b"11000000000000101000111101011100"), -- -7.05 + 5.01 = -2.04
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100101110000101000111101", b"00111111110101110000101001000000"), -- 6.4 + -4.72 = 1.68
	(b"01000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000001000000101011100001010010", b"11000000100010010100011110101110"), -- 3.88 + -8.17 = -4.29
	(b"11000001000001101000111101011100", b"00000000000000000000000000000000"),
	(b"01000001000001100011110101110001", b"10111100101000111101011000000000"), -- -8.41 + 8.39 = -0.0199995
	(b"11000000101111111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010110100011110101110001", b"11000001000101100110011001100110"), -- -5.99 + -3.41 = -9.4
	(b"01000001000101110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000111110101000111101011100", b"00111111110100001010001111011000"), -- 9.46 + -7.83 = 1.63
	(b"01000000111010010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000110011110101110000101001", b"01000001010111000101000111101100"), -- 7.29 + 6.48 = 13.77
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000101011100001010001111", b"11000000010101011100001010001111"), -- -1 + -2.34 = -3.34
	(b"01000000100100010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000111110000101000111101100", b"11000000010011100001010001111100"), -- 4.54 + -7.76 = -3.22
	(b"01000001000101101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111000011110101110000101001", b"01000001000111111000010100011111"), -- 9.41 + 0.56 = 9.97
	(b"01000000110100001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000110000100011110101110001", b"00111110111010111000010100100000"), -- 6.53 + -6.07 = 0.46
	(b"01000001000110110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000111101110101110000101001", b"01000001100010111000010100011111"), -- 9.71 + 7.73 = 17.44
	(b"01000000101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000101100001010001111010111", b"10111110110011001100110011010000"), -- 5.12 + -5.52 = -0.4
	(b"11000001000100010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111101000111101011100001010", b"11000001001001011001100110011001"), -- -9.07 + -1.28 = -10.35
	(b"01000001000101000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000001100000000000000000000", b"01000000110100000101000111101100"), -- 9.26 + -2.75 = 6.51
	(b"10111111111111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000001000001100011110101110001", b"01000000110011001100110011001110"), -- -1.99 + 8.39 = 6.4
	(b"01000000100001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000000100011110101110000101001"), -- 4.22 + -8.7 = -4.48
	(b"01000001000010111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111000010100011110101110001", b"01000001000000110000101000111101"), -- 8.73 + -0.54 = 8.19
	(b"01000000110001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101010111000010100100", b"01000001011101111101011100001010"), -- 6.15 + 9.34 = 15.49
	(b"01000001000110100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"01000001001010000010100011110110"), -- 9.64 + 0.87 = 10.51
	(b"01000001000111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111011101011100001010010", b"01000001100010110100011110101110"), -- 9.95 + 7.46 = 17.41
	(b"11000000011011010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000100011000010100011110110", b"11000001000000010111000010100100"), -- -3.71 + -4.38 = -8.09
	(b"01000000100001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000001000110011100001010001111", b"11000000101011000111101011100001"), -- 4.22 + -9.61 = -5.39
	(b"01000000101011011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111100110101110000101001000", b"01000000110101000111101011100001"), -- 5.43 + 1.21 = 6.64
	(b"11000001000101000000000000000000", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"11000001000101000010100011110110"), -- -9.25 + -0.01 = -9.26
	(b"11000000110100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111100001111010111000010100", b"11000000111101011100001010001111"), -- -6.62 + -1.06 = -7.68
	(b"11000000100110010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000100100001010001111010111", b"11000001000101001111010111000010"), -- -4.79 + -4.52 = -9.31
	(b"11000001000000011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000100101011100001010001111", b"11000001010011001100110011001100"), -- -8.12 + -4.68 = -12.8
	(b"01000000101111010001111010111000", b"00000000000000000000000000000000"),
	(b"01000001000001101110000101001000", b"01000001011001010111000010100100"), -- 5.91 + 8.43 = 14.34
	(b"11000000111100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000001000001100001010001111011", b"00111111010111000010100011111000"), -- -7.52 + 8.38 = 0.86
	(b"11000000011101010001111010111000", b"00000000000000000000000000000000"),
	(b"11000001000101100001010001111011", b"11000001010100110101110000101001"), -- -3.83 + -9.38 = -13.21
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011010111000010100100", b"01000000111110011110101110000101"), -- 4.1 + 3.71 = 7.81
	(b"11000000001010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000101000011001100110011010", b"01000000000110101110000101001000"), -- -2.63 + 5.05 = 2.42
	(b"01000000111101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000001000101010100011110101110", b"10111111110011100001010001111100"), -- 7.72 + -9.33 = -1.61
	(b"11000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000001000100100001010001111011"), -- -2.93 + -6.2 = -9.13
	(b"11000001000111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000101111010111000010100100", b"11000001011111000010100011110110"), -- -9.84 + -5.92 = -15.76
	(b"01000000111111110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111111011001100110011001101", b"01000001000111010001111010111000"), -- 7.97 + 1.85 = 9.82
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000111100011001100110011010", b"11000000111101100001010001111011"), -- -0.14 + -7.55 = -7.69
	(b"01000000100000001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000100000111101011100001010", b"01000001000000100110011001100110"), -- 4.03 + 4.12 = 8.15
	(b"11000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000000101011100001010001111", b"11000000100110110011001100110011"), -- -2.51 + -2.34 = -4.85
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110111000111101011100001", b"11000000010001011100001010001111"), -- 3.8 + -6.89 = -3.09
	(b"11000001000100010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000101000000101000111101100", b"11000001011000011001100110011010"), -- -9.09 + -5.01 = -14.1
	(b"11000000110000111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000101000101000111101011100", b"10111111100000111101011100001100"), -- -6.11 + 5.08 = -1.03
	(b"11000000100111100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"11000000010111000010100011110110"), -- -4.94 + 1.5 = -3.44
	(b"01000001000101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000100001000111101011100001", b"01000000101010011001100110011001"), -- 9.44 + -4.14 = 5.3
	(b"01000001000111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000001000111000010100011110110", b"01000001100111011100001010010000"), -- 9.96 + 9.76 = 19.72
	(b"01000000110111000111101011100001", b"00000000000000000000000000000000"),
	(b"11000001000100110000101000111101", b"11000000000100110011001100110010"), -- 6.89 + -9.19 = -2.3
	(b"11000001000100000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"11000001000000001010001111010111"), -- -9.03 + 0.99 = -8.04
	(b"11000000011101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000100000001010001111010111", b"11000000111111000010100011110110"), -- -3.86 + -4.02 = -7.88
	(b"01000000000011010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000011110100011110101110001", b"01000000110000111101011100001010"), -- 2.21 + 3.91 = 6.12
	(b"11000001000111101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001000010110000101000111101", b"11000001100101001111010111000010"), -- -9.93 + -8.69 = -18.62
	(b"01000000110101111010111000010100", b"00000000000000000000000000000000"),
	(b"11000001000111111101011100001010", b"11000000010100000000000000000000"), -- 6.74 + -9.99 = -3.25
	(b"01000001000010110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110010101110000101000111101", b"01000001000011101011100001010010"), -- 8.71 + 0.21 = 8.92
	(b"11000000110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111111011110101110000101001", b"11000001000001101110000101001000"), -- -6.56 + -1.87 = -8.43
	(b"11000000100101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000001000110101000111101011100", b"11000001011001001100110011001100"), -- -4.64 + -9.66 = -14.3
	(b"01000000000000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000111010111101011100001010", b"11000000101010111000010100011110"), -- 2.01 + -7.37 = -5.36
	(b"10111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000001000101001111010111000011", b"01000001000010111010111000010101"), -- -0.58 + 9.31 = 8.73
	(b"00111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"00111110011010111000010100100000"), -- 0.49 + -0.26 = 0.23
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001000010100011110110", b"01000001011011000010100011110110"), -- 6.5 + 8.26 = 14.76
	(b"01000001000010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001010000101000111101100", b"01000001001101000111101011100001"), -- 8.65 + 2.63 = 11.28
	(b"11000000101110010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111000111000010100011110110", b"11000000101001011100001010001111"), -- -5.79 + 0.61 = -5.18
	(b"10111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111010111000010100011110110", b"00111111000001010001111010111000"), -- -0.34 + 0.86 = 0.52
	(b"11000000111111111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111100110101110000101001000", b"11000000110110001111010111000010"), -- -7.99 + 1.21 = -6.78
	(b"10111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000100100111000010100011111", b"01000000100010001111010111000011"), -- -0.33 + 4.61 = 4.28
	(b"01000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001000110001111010111000011", b"11000000111001000111101011100010"), -- 2.42 + -9.56 = -7.14
	(b"11000000011000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000110011110101110000101001", b"01000000001111000010100011110110"), -- -3.54 + 6.48 = 2.94
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001000101100110011001100110"), -- -1.5 + -7.9 = -9.4
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"01000000101111000111101011100010"), -- 6.8 + -0.91 = 5.89
	(b"11000000110011010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"11000000101101111010111000010100"), -- -6.41 + 0.67 = -5.74
	(b"01000001000010010100011110101110", b"00000000000000000000000000000000"),
	(b"11000001000100000101000111101100", b"10111110111000010100011111000000"), -- 8.58 + -9.02 = -0.440001
	(b"11000000101001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000110010010100011110101110", b"00111111100100001010001111011000"), -- -5.16 + 6.29 = 1.13
	(b"01000000010100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101001000111101011100001", b"10111111111100011110101110000100"), -- 3.25 + -5.14 = -1.89
	(b"01000000101001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010100011110101110001", b"11000000010111110101110000101010"), -- 5.15 + -8.64 = -3.49
	(b"11000001000110000010100011110110", b"00000000000000000000000000000000"),
	(b"01000001000110001100110011001101", b"00111101001000111101011100000000"), -- -9.51 + 9.55 = 0.04
	(b"01000000100000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000100111011100001010001111", b"10111111010110011001100110011000"), -- 4.08 + -4.93 = -0.85
	(b"11000000101101000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000100011100110011001100110", b"11000001001000010100011110101110"), -- -5.63 + -4.45 = -10.08
	(b"01000001000010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000111010101110000101001000", b"01000001100000000111101011100010"), -- 8.72 + 7.34 = 16.06
	(b"01000000101110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000000010010001111010111000000"), -- 5.76 + -8.9 = -3.14
	(b"11000000111000000101000111101100", b"00000000000000000000000000000000"),
	(b"01000001000100000111101011100001", b"01000000000000010100011110101100"), -- -7.01 + 9.03 = 2.02
	(b"01000001000100000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000100100011001100110011010", b"01000000100011101011100001010010"), -- 9.01 + -4.55 = 4.46
	(b"10111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000000000001010001111010111", b"00111111101110000101000111101100"), -- -0.57 + 2.01 = 1.44
	(b"00111111111101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000001000001000111101011100001", b"01000001001000110000101000111101"), -- 1.91 + 8.28 = 10.19
	(b"11000000101001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100010100011110101110", b"11000000000110000101000111101100"), -- -5.15 + 2.77 = -2.38
	(b"11000000110101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000100001111010111000010100", b"11000000000111000010100011110110"), -- -6.68 + 4.24 = -2.44
	(b"11000000000111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000111011110000101000111101", b"01000000101000000101000111101011"), -- -2.46 + 7.47 = 5.01
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111110101111010111000010100101"), -- -0.42 + 0.79 = 0.37
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000111111111010111000010100", b"01000000111010100011110101110000"), -- -0.67 + 7.99 = 7.32
	(b"01000000111110010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111100101011100001010001111", b"01000001000011110101110000101001"), -- 7.79 + 1.17 = 8.96
	(b"00111111100001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110111000010100011110101110", b"00111111101111101011100001010010"), -- 1.05 + 0.44 = 1.49
	(b"11000000110000011110101110000101", b"00000000000000000000000000000000"),
	(b"11000001000000011110101110000101", b"11000001011000101110000101001000"), -- -6.06 + -8.12 = -14.18
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110100000000000000000000000"), -- -0.15 + 0.4 = 0.25
	(b"01000001000000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000101010010100011110101110", b"01000000001100101000111101011100"), -- 8.08 + -5.29 = 2.79
	(b"00111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111100000101000111101011100", b"00111111100011001100110011001101"), -- 0.08 + 1.02 = 1.1
	(b"01000000110011101011100001010010", b"00000000000000000000000000000000"),
	(b"11000001000000110101110000101001", b"10111111111000000000000000000000"), -- 6.46 + -8.21 = -1.75
	(b"11000000010111100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111110010001111010111000011"), -- -3.47 + 1.9 = -1.57
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111110001111010111000011", b"10111111011110101110000101001000"), -- 6.8 + -7.78 = -0.98
	(b"10111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000000101100001010001111010111"), -- -0.98 + 6.5 = 5.52
	(b"01000001000000100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011110101110000101001", b"01000001000111000101000111101011"), -- 8.15 + 1.62 = 9.77
	(b"11000001000011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101000000000000000000", b"11000001100100011001100110011010"), -- -8.95 + -9.25 = -18.2
	(b"01000000101100001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000100011110000101000111101", b"01000001001000000000000000000000"), -- 5.53 + 4.47 = 10
	(b"01000000100010101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"01000000100100001111010111000011"), -- 4.34 + 0.19 = 4.53
	(b"10111111110010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111101001010001111010111000", b"11000000001110000101000111101100"), -- -1.59 + -1.29 = -2.88
	(b"11000000110110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000001000000001100110011001101", b"11000001011011100011110101110001"), -- -6.84 + -8.05 = -14.89
	(b"01000001000101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111111000010100011110101110", b"01000000111101011100001010001110"), -- 9.44 + -1.76 = 7.68
	(b"10111111101011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000110000100011110101110001", b"11000000111011011100001010010000"), -- -1.36 + -6.07 = -7.43
	(b"11000001000011101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000100100010100011110101110", b"11000001010101110011001100110011"), -- -8.91 + -4.54 = -13.45
	(b"01000001000000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000100001010001111010111000", b"01000000011110101110000101001000"), -- 8.08 + -4.16 = 3.92
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001101110000101000111101", b"11000001001011110101110000101001"), -- -8.1 + -2.86 = -10.96
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101000010100011110110", b"10111110100010100011110101110000"), -- -6.9 + 6.63 = -0.27
	(b"01000000101100101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000001000111101011100001010", b"01000001000000100110011001100110"), -- 5.59 + 2.56 = 8.15
	(b"01000000001101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000101011100110011001100110", b"11000000001001011100001010001111"), -- 2.86 + -5.45 = -2.59
	(b"11000000001001011100001010001111", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000001001111001010001111010111"), -- -2.59 + -9.2 = -11.79
	(b"11000000101100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010110100011110101110001", b"11000001000011101110000101001000"), -- -5.52 + -3.41 = -8.93
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000111011000111101011100001", b"01000000110100011110101110000101"), -- -0.83 + 7.39 = 6.56
	(b"01000001000001001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000010010100011110101110001", b"01000001001101111000010100011111"), -- 8.31 + 3.16 = 11.47
	(b"01000000100110000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"01000000100001000111101011100001"), -- 4.75 + -0.61 = 4.14
	(b"11000001000101010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000100011111010111000010100", b"11000000100110101110000101001000"), -- -9.33 + 4.49 = -4.84
	(b"11000001000000100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000100111000111101011100001", b"11000001010100000111101011100010"), -- -8.14 + -4.89 = -13.03
	(b"01000000100010101110000101001000", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"01000000100010001111010111000011"), -- 4.34 + -0.06 = 4.28
	(b"11000000110011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000001000101011001100110011010", b"01000000001101111010111000010110"), -- -6.48 + 9.35 = 2.87
	(b"01000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000111101010001111010111000", b"01000001001010100001010001111011"), -- 2.97 + 7.66 = 10.63
	(b"01000000101011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000001000001000111101011100001", b"01000001010111000010100011110110"), -- 5.48 + 8.28 = 13.76
	(b"11000000010011101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000000010111000010100011111", b"11000000101011010001111010111000"), -- -3.23 + -2.18 = -5.41
	(b"01000000010101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110001010001111010111000", b"11000000001100111101011100001010"), -- 3.35 + -6.16 = -2.81
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101010001111010111000011", b"11000000101111000010100011110110"), -- -0.6 + -5.28 = -5.88
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100001111010111000010100", b"11000000110010111000010100011111"), -- -5.3 + -1.06 = -6.36
	(b"01000000111000001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"01000000110011101011100001010010"), -- 7.03 + -0.57 = 6.46
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000100110000000000000000000", b"01000000100000111000010100011111"), -- -0.64 + 4.75 = 4.11
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001010001111010111000", b"01000000000110100011110101110000"), -- 4.2 + -1.79 = 2.41
	(b"11000000110111100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101010111000010100011111", b"11000001000001001010001111010111"), -- -6.95 + -1.34 = -8.29
	(b"11000000110101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110001000111101011100001", b"10111111000000101000111101100000"), -- -6.65 + 6.14 = -0.51
	(b"01000001000001100011110101110001", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000001100001110001111010111000"), -- 8.39 + 8.5 = 16.89
	(b"11000000111001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000111010001111010111000", b"01000000001010101110000101000110"), -- -7.15 + 9.82 = 2.67
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100111000010100011111", b"01000001010101101000111101011100"), -- 8.8 + 4.61 = 13.41
	(b"11000000101100100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"11000000100111010111000010100100"), -- -5.57 + 0.65 = -4.92
	(b"11000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111111101011100001010001111", b"11000000101010101110000101001000"), -- -3.42 + -1.92 = -5.34
	(b"10111111110110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000101011010111000010100100", b"11000000111001000010100011110110"), -- -1.71 + -5.42 = -7.13
	(b"01000000111000101110000101001000", b"00000000000000000000000000000000"),
	(b"01000001000101001111010111000011", b"01000001100000110011001100110100"), -- 7.09 + 9.31 = 16.4
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010000111101011100001", b"11000000100001000010100011110101"), -- 4.4 + -8.53 = -4.13
	(b"11000001000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111101101011100001010001111", b"11000001000110010100011110101110"), -- -8.16 + -1.42 = -9.58
	(b"11000001000110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000001010001110011001100110011"), -- -9.65 + -2.8 = -12.45
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001010010000000000000000000"), -- -2.8 + -9.7 = -12.5
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011111100001010001111011", b"01000001000011000101000111101100"), -- 4.8 + 3.97 = 8.77
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000000001011100001010001111", b"10111111101001100110011001100110"), -- 0.79 + -2.09 = -1.3
	(b"11000000100101111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000010101111010111000010100", b"10111111101011110101110000101000"), -- -4.74 + 3.37 = -1.37
	(b"11000000110110101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000111111111010111000010100", b"00111111100101000111101011100000"), -- -6.83 + 7.99 = 1.16
	(b"11000000101001001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101110011001100110011010", b"11000000110100110011001100110100"), -- -5.15 + -1.45 = -6.6
	(b"01000000001100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000110001110101110000101001", b"11000000010111100001010001111011"), -- 2.76 + -6.23 = -3.47
	(b"10111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111101111010111000010100100", b"00111111101101000111101011100001"), -- -0.07 + 1.48 = 1.41
	(b"01000000011100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100110110011001100110011", b"01000001000010011001100110011010"), -- 3.75 + 4.85 = 8.6
	(b"00111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000100011110000101000111101"), -- 0.87 + 3.6 = 4.47
	(b"01000000111110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000110010001111010111000011", b"01000001011000011110101110000110"), -- 7.84 + 6.28 = 14.12
	(b"11000000010011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000001000001101110000101001000", b"11000001001110101011100001010010"), -- -3.24 + -8.43 = -11.67
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000001000010011110101110000101", b"01000000111110101000111101011100"), -- -0.79 + 8.62 = 7.83
	(b"01000001000000101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000001010000101000111101100", b"01000000101100010100011110101110"), -- 8.17 + -2.63 = 5.54
	(b"11000001000100001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"11000001000000001111010111000011"), -- -9.05 + 0.99 = -8.06
	(b"11000001000010011110101110000101", b"00000000000000000000000000000000"),
	(b"11000001000101001111010111000011", b"11000001100011110111000010100100"), -- -8.62 + -9.31 = -17.93
	(b"01000001000111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000100101000111101011100001", b"01000000101000111101011100001011"), -- 9.76 + -4.64 = 5.12
	(b"01000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000111001110000101000111101", b"11000000010101011100001010001110"), -- 3.88 + -7.22 = -3.34
	(b"10111111100001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000111100010100011110101110", b"01000000110011110101110000101001"), -- -1.06 + 7.54 = 6.48
	(b"11000000101101111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000010000011110101110000101", b"11000000001011010111000010100011"), -- -5.74 + 3.03 = -2.71
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000001000001001111010111000011", b"11000000111100001010001111011000"), -- 0.79 + -8.31 = -7.52
	(b"01000001000111011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000111111000010100011110110", b"00111111111111010111000010100000"), -- 9.86 + -7.88 = 1.98
	(b"01000000010001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000101101101011100001010010", b"11000000001010000101000111101100"), -- 3.08 + -5.71 = -2.63
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100010100011110101110", b"11000001000001000101000111101100"), -- -6 + -2.27 = -8.27
	(b"10111111110110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111111011000111101011100001011"), -- -1.69 + 0.8 = -0.89
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000001111100001010001111011", b"01000000000100000000000000000000"), -- -0.72 + 2.97 = 2.25
	(b"11000000101001000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000100110111000010100011111", b"11000001000111111101011100001010"), -- -5.13 + -4.86 = -9.99
	(b"01000000010100011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000100000000101000111101100", b"01000000111010010100011110101110"), -- 3.28 + 4.01 = 7.29
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000100010100011110101110001", b"01000000011000101000111101011101"), -- -0.78 + 4.32 = 3.54
	(b"11000000110111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000010110001111010111000011", b"11000001001001001111010111000011"), -- -6.92 + -3.39 = -10.31
	(b"10111111110010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000010010101110000101001000", b"11000000100101111010111000010101"), -- -1.57 + -3.17 = -4.74
	(b"11000000110100010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000011100000000000000000000", b"11000001001001001010001111010111"), -- -6.54 + -3.75 = -10.29
	(b"01000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101100000101000111101100", b"01000001010000011100001010010000"), -- 6.6 + 5.51 = 12.11
	(b"01000001000000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010001010001111010111000", b"01000000101000100011110101110000"), -- 8.15 + -3.08 = 5.07
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000101111010001111010111000", b"11000000101101010111000010100100"), -- 0.24 + -5.91 = -5.67
	(b"01000001000010101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000010101110000101000111101", b"01000000101010011110101110000110"), -- 8.67 + -3.36 = 5.31
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000011100111101011100001010", b"01000000010001011100001010001111"), -- -0.72 + 3.81 = 3.09
	(b"01000000110001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010101100110011001100110", b"01000001000110000000000000000000"), -- 6.15 + 3.35 = 9.5
	(b"00111111101101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111100010100011110101110001", b"01000000000111110101110000101001"), -- 1.41 + 1.08 = 2.49
	(b"01000000001001000111101011100001", b"00000000000000000000000000000000"),
	(b"01000001000100110101110000101001", b"01000001001111000111101011100001"), -- 2.57 + 9.21 = 11.78
	(b"11000000011000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000000111101000111101011100001"), -- -3.54 + -4.1 = -7.64
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111101010001111010111000", b"01000000101001010001111010111000"), -- -2.5 + 7.66 = 5.16
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000001000000000101000111101100", b"11000001000011001100110011001101"), -- -0.78 + -8.02 = -8.8
	(b"11000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110101000111101011100001010", b"11000000010001100110011001100111"), -- -3.42 + 0.32 = -3.1
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111100100011110101110000101", b"10111111100011110101110000101001"), -- 0.02 + -1.14 = -1.12
	(b"01000000111111111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111110010100011110101110001", b"01000001000110010001111010111000"), -- 7.99 + 1.58 = 9.57
	(b"10111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000110011110101110000101001", b"11000000110100000000000000000000"), -- -0.02 + -6.48 = -6.5
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100111101011100001010", b"01000001000111101011100001010010"), -- 3.3 + 6.62 = 9.92
	(b"10111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000010000011110101110000101", b"00111111101111000010100011110110"), -- -1.56 + 3.03 = 1.47
	(b"01000000101000001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000100110101000111101011100", b"00111110010011001100110011100000"), -- 5.03 + -4.83 = 0.2
	(b"01000001000001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000001000000101011100001010010", b"01000001100000111110101110000101"), -- 8.32 + 8.17 = 16.49
	(b"11000001000100101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000110100001111010111000011", b"11000001011110110000101000111110"), -- -9.16 + -6.53 = -15.69
	(b"01000000010000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000110101010111000010100100", b"01000001000110110101110000101001"), -- 3.04 + 6.67 = 9.71
	(b"11000000101101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111101011001100110011001101", b"11000000111000100011110101110000"), -- -5.72 + -1.35 = -7.07
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100011110101110000101", b"10111111101010111000010100100000"), -- -5.9 + 4.56 = -1.34
	(b"11000000011011000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000101100001111010111000011", b"11000001000100111000010100011111"), -- -3.69 + -5.53 = -9.22
	(b"11000000000011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000101111101011100001010010", b"01000000011011110101110000101001"), -- -2.22 + 5.96 = 3.74
	(b"01000000100110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000101111110101110000101001", b"10111111100100011110101110000100"), -- 4.84 + -5.98 = -1.14
	(b"01000000110000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000100111011100001010001111", b"00111111100110000101000111101100"), -- 6.12 + -4.93 = 1.19
	(b"11000001000011010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000110000100011110101110001", b"11000000001011111111111111111110"), -- -8.82 + 6.07 = -2.75
	(b"11000000010100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000110010111000010100011111", b"01000000010000110011001100110100"), -- -3.31 + 6.36 = 3.05
	(b"01000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000110000010100011110101110", b"01000001001000000101000111101100"), -- 3.98 + 6.04 = 10.02
	(b"11000000101011000010100011110110", b"00000000000000000000000000000000"),
	(b"01000001000010001111010111000011", b"01000000010010111000010100100000"), -- -5.38 + 8.56 = 3.18
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110010001111010111000011", b"10111111101010100011110101110001"), -- -2.9 + 1.57 = -1.33
	(b"00111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000110100111000010100011111", b"01000000110110111101011100001010"), -- 0.26 + 6.61 = 6.87
	(b"11000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000001000100010111000010100100", b"11000001010000001111010111000011"), -- -2.97 + -9.09 = -12.06
	(b"11000000110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111110101110000101000111101", b"11000001000000111101011100001010"), -- -6.56 + -1.68 = -8.24
	(b"10111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110100011110101110000101", b"10111111000010100011110101110000"), -- -0.95 + 0.41 = -0.54
	(b"01000000011111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100111000010100011110110", b"10111111011011100001010001111100"), -- 3.95 + -4.88 = -0.93
	(b"00111111101010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000101101010001111010111000", b"01000000110111111010111000010100"), -- 1.33 + 5.66 = 6.99
	(b"11000000101101100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"11000000101111100110011001100110"), -- -5.69 + -0.26 = -5.95
	(b"11000001000110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"11000001000011100011110101110001"), -- -9.68 + 0.79 = -8.89
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100010001010001111010111", b"11000001000000101011100001010010"), -- -3.9 + -4.27 = -8.17
	(b"10111111100100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111111001111010111000010100", b"00111111001011100001010001111010"), -- -1.13 + 1.81 = 0.68
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100100100011110101110001", b"01000000101100100011110101110001"), -- 1 + 4.57 = 5.57
	(b"11000001000010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001111010111000010100", b"11000000100111011100001010010000"), -- -8.55 + 3.62 = -4.93
	(b"10111111111010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000111010111000010100011111", b"11000001000100110011001100110011"), -- -1.84 + -7.36 = -9.2
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000010101110000101001000", b"00111111011011100001010001111000"), -- 3.1 + -2.17 = 0.93
	(b"11000000000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110100001010001111011", b"11000001001111111010111000010100"), -- -2.35 + -9.63 = -11.98
	(b"11000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000110000111101011100001010", b"11000001000011110000101000111101"), -- -2.82 + -6.12 = -8.94
	(b"01000001000101111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"01000001001000011110101110000101"), -- 9.48 + 0.64 = 10.12
	(b"11000000111101110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000110001100001010001111011", b"11000001010111101011100001010010"), -- -7.73 + -6.19 = -13.92
	(b"10111111100010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000100011010001111010111000", b"11000000101011111010111000010100"), -- -1.08 + -4.41 = -5.49
	(b"00111111011011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000001000001010100011110101110", b"01000001000101000010100011110110"), -- 0.93 + 8.33 = 9.26
	(b"11000000110010111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000011100101000111101011100", b"11000001001000101000111101011100"), -- -6.37 + -3.79 = -10.16
	(b"11000000100100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110110100011110101110001", b"01000000000100010100011110101110"), -- -4.55 + 6.82 = 2.27
	(b"11000000111011000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000010111110101110000101001", b"11000001001011100001010001111011"), -- -7.39 + -3.49 = -10.88
	(b"01000000110110100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111110001111010111000010100", b"01000001000001100001010001111011"), -- 6.82 + 1.56 = 8.38
	(b"11000001000011000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"11000001000001010001111010111000"), -- -8.75 + 0.43 = -8.32
	(b"01000001000011001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001011111111101011100001010"), -- 8.79 + 7.2 = 15.99
	(b"01000000001111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000001000001000101000111101100", b"01000001001101000010100011110110"), -- 2.99 + 8.27 = 11.26
	(b"11000001000001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100110001010001111010111", b"11000001010100011110101110000110"), -- -8.35 + -4.77 = -13.12
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110111010111000010100", b"11000000101010101000111101011011"), -- 4.4 + -9.73 = -5.33
	(b"11000000101011110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111110100011110101110000101", b"11000000111000111000010100011110"), -- -5.47 + -1.64 = -7.11
	(b"01000000010100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000111101011100001010001111", b"01000001001011111101011100001010"), -- 3.31 + 7.68 = 10.99
	(b"01000001000101001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000010100111101011100001010", b"01000001010010011001100110011010"), -- 9.29 + 3.31 = 12.6
	(b"00111111110101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000000001101000111101011100010"), -- 1.68 + -4.5 = -2.82
	(b"11000000111100010100011110101110", b"00000000000000000000000000000000"),
	(b"01000001000011001010001111010111", b"00111111101000000000000000000000"), -- -7.54 + 8.79 = 1.25
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000001100001010001111010111", b"11000000010010000101000111101100"), -- -0.37 + -2.76 = -3.13
	(b"11000000000001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000101101000010100011110110", b"11000000111101111010111000010100"), -- -2.11 + -5.63 = -7.74
	(b"11000001000100101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000100101000111101011100001", b"11000000100100001010001111010111"), -- -9.16 + 4.64 = -4.52
	(b"11000000101101100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000011010101110000101001000", b"11000000000000010100011110101110"), -- -5.69 + 3.67 = -2.02
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000010111000010100011111", b"00111101101000111101011100100000"), -- -2.1 + 2.18 = 0.0800002
	(b"01000000100000000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000101100011001100110011010", b"01000001000110001111010111000011"), -- 4.01 + 5.55 = 9.56
	(b"11000000101000000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000011011010111000010100100", b"11000001000010111000010100011111"), -- -5.01 + -3.71 = -8.72
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000010101110000101001000", b"00111111000101000111101011100000"), -- -8.1 + 8.68 = 0.58
	(b"01000000111000001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111100011110101110000101001", b"01000000101111010001111010111001"), -- 7.03 + -1.12 = 5.91
	(b"10111111111111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111111101110000101000111101", b"10111101001000111101011100100000"), -- -1.97 + 1.93 = -0.0400001
	(b"01000000111101111010111000010100", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"01000000111101100001010001111010"), -- 7.74 + -0.05 = 7.69
	(b"11000000110100100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010000001010001111010111", b"11000000011000111101011100001011"), -- -6.57 + 3.01 = -3.56
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010110000101000111101", b"00111111001100001010001111010000"), -- -8 + 8.69 = 0.69
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011101011100001010010", b"01000000100111011100001010010000"), -- 2.2 + 2.73 = 4.93
	(b"10111111101000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111110011100001010001111011", b"00111110101011100001010001111100"), -- -1.27 + 1.61 = 0.34
	(b"01000000101110100011110101110001", b"00000000000000000000000000000000"),
	(b"01000001000010111000010100011111", b"01000001011010001010001111011000"), -- 5.82 + 8.72 = 14.54
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000101100110011001100110", b"01000001010000001100110011001100"), -- 9.7 + 2.35 = 12.05
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100011111010111000010100", b"11000000010011010111000010100100"), -- -7.7 + 4.49 = -3.21
	(b"01000001000110010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000000101100110011001100110", b"01000001001111101011100001010010"), -- 9.57 + 2.35 = 11.92
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000100000111000010100011111", b"11000000011110001111010111000011"), -- 0.22 + -4.11 = -3.89
	(b"01000001000101101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000100010000101000111101100", b"01000001010110110000101000111110"), -- 9.43 + 4.26 = 13.69
	(b"01000000111001000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000001101111010111000010100", b"01000000100010000101000111101100"), -- 7.13 + -2.87 = 4.26
	(b"00111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000010100000000000000000000", b"11000000001101011100001010001111"), -- 0.41 + -3.25 = -2.84
	(b"11000001000110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001110011001100110011", b"11000001100100000000000000000000"), -- -9.55 + -8.45 = -18
	(b"01000000110101101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000101000100011110101110001", b"00111111110100011110101110000100"), -- 6.71 + -5.07 = 1.64
	(b"11000000100011011100001010001111", b"00000000000000000000000000000000"),
	(b"11000001000000101000111101011100", b"11000001010010010111000010100100"), -- -4.43 + -8.16 = -12.59
	(b"01000000100000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000001000110001100110011001101", b"01000001010110010111000010100100"), -- 4.04 + 9.55 = 13.59
	(b"01000000100101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000011100101000111101011100", b"00111111011000111101011100001000"), -- 4.68 + -3.79 = 0.89
	(b"00111111100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000001111010111000011", b"11000000110111010001111010111001"), -- 1.15 + -8.06 = -6.91
	(b"01000000111010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"01000000110100100011110101110001"), -- 7.36 + -0.79 = 6.57
	(b"10111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000011000010100011110101110", b"01000000001100011110101110000101"), -- -0.74 + 3.52 = 2.78
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101001100001010001111011", b"01000001011100010111000010100100"), -- 9.9 + 5.19 = 15.09
	(b"11000000100110111101011100001010", b"00000000000000000000000000000000"),
	(b"01000001000101011001100110011010", b"01000000100011110101110000101010"), -- -4.87 + 9.35 = 4.48
	(b"00111111100100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"01000000000001000111101011100001"), -- 1.13 + 0.94 = 2.07
	(b"10111111101000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111110100001010001111010111", b"11000000001110001111010111000010"), -- -1.26 + -1.63 = -2.89
	(b"11000001000101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011011001100110011010", b"11000001100100100110011001100110"), -- -9.45 + -8.85 = -18.3
	(b"01000000110010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000101101101011100001010010", b"01000001010000001100110011001101"), -- 6.34 + 5.71 = 12.05
	(b"10111111111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111111010001111010111000", b"01000000101111101011100001010010"), -- -1.95 + 7.91 = 5.96
	(b"11000000111010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011010001111010111000011", b"11000001001011100011110101110001"), -- -7.25 + -3.64 = -10.89
	(b"00111111100111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111100001111010111000010100", b"01000000000100110011001100110011"), -- 1.24 + 1.06 = 2.3
	(b"10111111110010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000010000101000111101011100", b"11000000100100111000010100011111"), -- -1.57 + -3.04 = -4.61
	(b"01000001000000011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"01000000111111100001010001111010"), -- 8.11 + -0.17 = 7.94
	(b"10111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000011101000111101011100001", b"01000000010111110101110000101001"), -- -0.33 + 3.82 = 3.49
	(b"11000000101101100001010001111011", b"00000000000000000000000000000000"),
	(b"11000001000001010100011110101110", b"11000001011000000101000111101100"), -- -5.69 + -8.33 = -14.02
	(b"11000000111000000101000111101100", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"11000000111000011110101110000110"), -- -7.01 + -0.05 = -7.06
	(b"11000001000010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100110111000010100011111", b"11000000011011000010100011110110"), -- -8.55 + 4.86 = -3.69
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000001000010100110011001100110", b"01000001000101000101000111101011"), -- 0.62 + 8.65 = 9.27
	(b"11000000101010101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"11000000110000111101011100001010"), -- -5.34 + -0.78 = -6.12
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001010111000010100011111", b"01000000001010111000010100011111"), -- 0 + 2.68 = 2.68
	(b"11000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000001000111100011110101110001", b"01000000101111010001111010111001"), -- -3.98 + 9.89 = 5.91
	(b"11000000000011101011100001010010", b"00000000000000000000000000000000"),
	(b"11000001000111010001111010111000", b"11000001010000001100110011001100"), -- -2.23 + -9.82 = -12.05
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100110000101000111101", b"01000001000110010111000010100011"), -- 0.4 + 9.19 = 9.59
	(b"11000001000001110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000011100001010001111010111", b"11000001010000111000010100011111"), -- -8.46 + -3.76 = -12.22
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000100011110101110000101", b"10111111101010100011110101110000"), -- -1.9 + 0.57 = -1.33
	(b"11000001000011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000101011011100001010001111", b"11000001011001100011110101110000"), -- -8.96 + -5.43 = -14.39
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001011100001010001111", b"00111110010000101000111101011000"), -- -1.9 + 2.09 = 0.19
	(b"01000000101110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111111101011100001010010", b"11000000000011010111000010100100"), -- 5.75 + -7.96 = -2.21
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100000111000010100011111", b"01000000111000000101000111101100"), -- 2.9 + 4.11 = 7.01
	(b"10111111101101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000010000010100011110101110", b"00111111110011001100110011001101"), -- -1.42 + 3.02 = 1.6
	(b"01000000000100101000111101011100", b"00000000000000000000000000000000"),
	(b"11000001000011010001111010111000", b"11000000110100001111010111000010"), -- 2.29 + -8.82 = -6.53
	(b"01000001000000100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000101100010100011110101110", b"01000000001001100110011001101000"), -- 8.14 + -5.54 = 2.6
	(b"00111111101111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000100111100001010001111011", b"11000000010111010111000010100100"), -- 1.48 + -4.94 = -3.46
	(b"11000000010110100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000111000010100011110101110", b"11000001001001110011001100110011"), -- -3.41 + -7.04 = -10.45
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"01000000010110011001100110011000"), -- 9.7 + -6.3 = 3.4
	(b"01000001000001110101110000101001", b"00000000000000000000000000000000"),
	(b"01000001000111001111010111000011", b"01000001100100100010100011110110"), -- 8.46 + 9.81 = 18.27
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000110001110101110000101001", b"11000000110101010001111010111000"), -- -0.43 + -6.23 = -6.66
	(b"11000000011100111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111110010100011110101110001", b"11000000000011101011100001010010"), -- -3.81 + 1.58 = -2.23
	(b"01000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000101110001010001111010111", b"11000000001100110011001100110011"), -- 2.97 + -5.77 = -2.8
	(b"11000000000000001010001111010111", b"00000000000000000000000000000000"),
	(b"01000001000000111010111000010100", b"01000000110001110000101000111100"), -- -2.01 + 8.23 = 6.22
	(b"11000000110100111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"11000000111001011100001010010000"), -- -6.61 + -0.57 = -7.18
	(b"01000000110010011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000001111100001010001111011", b"01000001000101000111101011100001"), -- 6.31 + 2.97 = 9.28
	(b"11000000000101010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000110110101000111101011100", b"11000001000100101000111101011100"), -- -2.33 + -6.83 = -9.16
	(b"01000000101010110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000011110101110000101001", b"01000000100110010100011110101110"), -- 5.35 + -0.56 = 4.79
	(b"01000001000110111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000100010111000010100011111", b"01000000101010111101011100001001"), -- 9.73 + -4.36 = 5.37
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110011110101110000101001", b"11000000101010001111010111000010"), -- 1.2 + -6.48 = -5.28
	(b"11000000110110111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111000111000010100011110110", b"11000000110010000101000111101011"), -- -6.87 + 0.61 = -6.26
	(b"01000001000111100011110101110001", b"00000000000000000000000000000000"),
	(b"01000001000110000111101011100001", b"01000001100110110101110000101001"), -- 9.89 + 9.53 = 19.42
	(b"11000000100111011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000011001111010111000010100", b"10111111101001111010111000010100"), -- -4.93 + 3.62 = -1.31
	(b"11000000111000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"11000000000000010100011110101110"), -- -7.12 + 5.1 = -2.02
	(b"01000000111000111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000110000001111010111000011", b"00111111100010100011110101110000"), -- 7.11 + -6.03 = 1.08
	(b"11000000111101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000111011100110011001100110", b"10111110100010100011110101110000"), -- -7.72 + 7.45 = -0.27
	(b"01000001000011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000001000110010100011110101110", b"10111111000111101011100001010000"), -- 8.96 + -9.58 = -0.62
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"11000000101111110000101000111110"), -- -5.4 + -0.57 = -5.97
	(b"00111111111010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000101111100110011001100110", b"11000000100000111000010100011110"), -- 1.84 + -5.95 = -4.11
	(b"01000000101110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000100100111000010100011111", b"01000001001001110011001100110100"), -- 5.84 + 4.61 = 10.45
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000111111000010100011110110", b"11000000111101000111101011100010"), -- 0.24 + -7.88 = -7.64
	(b"01000000110100111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111111101110000101000111101", b"01000001000010001010001111010111"), -- 6.61 + 1.93 = 8.54
	(b"01000000101101111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000101001000111101011100001", b"01000001001011100001010001111010"), -- 5.74 + 5.14 = 10.88
	(b"11000000110011000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111111000000000000000000000", b"11000000100101000111101011100001"), -- -6.39 + 1.75 = -4.64
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001111010111000010100", b"01000001010001111010111000010100"), -- 4 + 8.48 = 12.48
	(b"11000000010000011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000000000011110101110000101"), -- -3.03 + 1 = -2.03
	(b"01000000110010111101011100001010", b"00000000000000000000000000000000"),
	(b"11000001000001101000111101011100", b"11000000000000101000111101011100"), -- 6.37 + -8.41 = -2.04
	(b"01000000001011010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000011111001100110011001101", b"01000000110101010001111010111000"), -- 2.71 + 3.95 = 6.66
	(b"01000000110111011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000101101011100001010001111", b"00111111101000000000000000000000"), -- 6.93 + -5.68 = 1.25
	(b"01000000101011111010111000010100", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000001011000110000101000111101"), -- 5.49 + 8.7 = 14.19
	(b"01000000110101101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000100101100001010001111011", b"01000000000000010100011110101110"), -- 6.71 + -4.69 = 2.02
	(b"11000000000010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"10111111101001111010111000010101"), -- -2.18 + 0.87 = -1.31
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101001110000101000111101", b"11000001001010000101000111101100"), -- -5.3 + -5.22 = -10.52
	(b"01000000110110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000100101001100110011001101", b"01000000000011000010100011110110"), -- 6.84 + -4.65 = 2.19
	(b"01000001000100111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000011011110101110000101001", b"01000000101011110101110000101010"), -- 9.22 + -3.74 = 5.48
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001101111010111000010100", b"11000001000111111000010100011110"), -- -7.1 + -2.87 = -9.97
	(b"11000000111011000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000111000000101000111101100", b"10111110110000101000111101010000"), -- -7.39 + 7.01 = -0.38
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110001110000101000111101", b"11000000011110101110000101000111"), -- 2.3 + -6.22 = -3.92
	(b"01000000100011010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000101010010100011110101110", b"01000001000110110011001100110011"), -- 4.41 + 5.29 = 9.7
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110011100110011001100110", b"01000000010101100110011001100110"), -- -3.1 + 6.45 = 3.35
	(b"01000000111001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"01000000111100001111010111000010"), -- 7.16 + 0.37 = 7.53
	(b"11000000011011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000001000011000101000111101100", b"11000001010001111101011100001011"), -- -3.72 + -8.77 = -12.49
	(b"01000000100111110000101000111101", b"00000000000000000000000000000000"),
	(b"01000001000001011110101110000101", b"01000001010101010111000010100100"), -- 4.97 + 8.37 = 13.34
	(b"01000001000001001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"01000000101001100001010001111011"), -- 8.29 + -3.1 = 5.19
	(b"11000000111111111010111000010100", b"00000000000000000000000000000000"),
	(b"01000001000101011100001010001111", b"00111111101011110101110000101000"), -- -7.99 + 9.36 = 1.37
	(b"01000001000100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110101110000101001000", b"01000000101101110101110000101000"), -- 9.15 + -3.42 = 5.73
	(b"01000000111010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000001000111100001010001111011", b"01000001100010011100001010010000"), -- 7.34 + 9.88 = 17.22
	(b"11000000001010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000110110110011001100110011", b"01000000100001011100001010001111"), -- -2.67 + 6.85 = 4.18
	(b"01000000100110111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000111010100011110101110001", b"11000000000111001100110011001110"), -- 4.87 + -7.32 = -2.45
	(b"01000001000001111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000011110101110000101001000", b"01000000100100011001100110011010"), -- 8.47 + -3.92 = 4.55
	(b"01000001000001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101000101000111101011100", b"01000000010010101110000101001000"), -- 8.25 + -5.08 = 3.17
	(b"11000000101000001111010111000011", b"00000000000000000000000000000000"),
	(b"01000001000100100001010001111011", b"01000000100000110011001100110011"), -- -5.03 + 9.13 = 4.1
	(b"00111111110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011101011100001010010", b"11000000000001010001111010111000"), -- 1.65 + -3.73 = -2.08
	(b"01000001000111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000001000101000111101011100", b"01000001010001101011100001010010"), -- 9.88 + 2.54 = 12.42
	(b"00111111100010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000111000111101011100001010", b"11000000110000001111010111000010"), -- 1.09 + -7.12 = -6.03
	(b"01000000100111000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110100101000111101011100001", b"01000000100100110011001100110011"), -- 4.89 + -0.29 = 4.6
	(b"01000001000011101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"01000000001101000111101011100010"), -- 8.92 + -6.1 = 2.82
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000010001111010111000010100", b"11000000011111000010100011110101"), -- -0.82 + -3.12 = -3.94
	(b"11000000111011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000000001000111101011100001", b"11000000101010111101011100001010"), -- -7.44 + 2.07 = -5.37
	(b"11000000100011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000101000010100011110101110", b"11000001000101111010111000010100"), -- -4.44 + -5.04 = -9.48
	(b"00111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000010100111101011100001010", b"11000000001101000111101011100001"), -- 0.49 + -3.31 = -2.82
	(b"01000000001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000100001101011100001010010", b"01000000110110001010001111010111"), -- 2.56 + 4.21 = 6.77

	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"10111111000111000010100011110110"), -- -0.14 + -0.47 = -0.61
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111101100011110101110000101001", b"10111110110111000010100011110110"), -- -0.36 + -0.07 = -0.43
	(b"00111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111001101011100001010001111", b"00111111010001010001111010111000"), -- 0.06 + 0.71 = 0.77
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111100110000101000111101100"), -- -0.39 + -0.8 = -1.19
	(b"10111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"10111110101111010111000010100100"), -- -0.33 + -0.04 = -0.37
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111001110000101000111101100"), -- -0.72 + -0 = -0.72
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111100001111010111000010101"), -- 0.6 + 0.46 = 1.06
	(b"00111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"00111111011101011100001010001111"), -- 0.71 + 0.25 = 0.96
	(b"10111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"10111110011101011100001010001111"), -- -0.08 + -0.16 = -0.24
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111011011100001010001111011", b"00111111101001111010111000010100"), -- 0.38 + 0.93 = 1.31
	(b"00111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"00111111011101011100001010010000"), -- 0.68 + 0.28 = 0.96
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"10111111101000010100011110101110"), -- -0.43 + -0.83 = -1.26
	(b"10111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"10111111110010111000010100011111"), -- -0.74 + -0.85 = -1.59
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"10111111100010111000010100011111"), -- -0.24 + -0.85 = -1.09
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"00111110101010001111010111000011"), -- 0.02 + 0.31 = 0.33
	(b"00111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110110100011110101110000101", b"00111111000001111010111000010100"), -- 0.12 + 0.41 = 0.53
	(b"00111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110000110011001100110011010", b"00111111010101000111101011100010"), -- 0.68 + 0.15 = 0.83
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111100101011100001010010000"), -- 0.63 + 0.54 = 1.17
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001010111000010100011111", b"10111111001110101110000101001000"), -- -0.06 + -0.67 = -0.73
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111010001010001111010111000", b"10111111110101000111101011100001"), -- -0.89 + -0.77 = -1.66
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111001110000101000111101100"), -- -0.42 + -0.3 = -0.72
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110000001010001111010111000", b"10111111000001010001111010111000"), -- -0.39 + -0.13 = -0.52
	(b"10111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001101011100001010001111", b"10111111100001111010111000010100"), -- -0.35 + -0.71 = -1.06
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111011001100110011001100110"), -- -0.37 + -0.53 = -0.9
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111110101110000101000111101100", b"00111111001000010100011110101110"), -- 0.27 + 0.36 = 0.63
	(b"00111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111110111101011100001010010"), -- 0.84 + 0.9 = 1.74
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111110010011001100110011001101"), -- -0.01 + -0.19 = -0.2
	(b"10111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"10111111101011100001010001111011"), -- -0.51 + -0.85 = -1.36
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111110100001010001111010111000", b"00111111000001111010111000010100"), -- 0.27 + 0.26 = 0.53
	(b"00111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111001000111101011100001010"), -- 0.18 + 0.46 = 0.64
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111001100001010001111010111", b"00111111100111010111000010100100"), -- 0.54 + 0.69 = 1.23
	(b"10111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111001011100001010001111011", b"10111111011100110011001100110100"), -- -0.27 + -0.68 = -0.95
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111100101011100001010001111"), -- -0.48 + -0.69 = -1.17
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101101110000101000111101100", b"10111110000011110101110000101001"), -- -0.05 + -0.09 = -0.14
	(b"00111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111110110000101000111101100"), -- 0.88 + 0.81 = 1.69
	(b"10111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111000010100011110101110001", b"10111111100101000111101011100010"), -- -0.62 + -0.54 = -1.16
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111110110101110000101001000"), -- -0.81 + -0.9 = -1.71
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111111010010100011110101110001"), -- 0.74 + 0.05 = 0.79
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"00111111101010111000010100011111"), -- 0.37 + 0.97 = 1.34
	(b"00111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"00111111010111000010100011110110"), -- 0.58 + 0.28 = 0.86
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111101111101011100001010001111", b"00111111001100001010001111010111"), -- 0.57 + 0.12 = 0.69
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111101100011110101110000101001", b"10111110101100110011001100110011"), -- -0.28 + -0.07 = -0.35
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111110110000101000111101011100"), -- 0.3 + 0.08 = 0.38
	(b"10111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"10111111011110000101000111101100"), -- -0.22 + -0.75 = -0.97
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111110101111010111000010100100"), -- 0.24 + 0.13 = 0.37
	(b"10111111011011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111101110000101000111101100"), -- -0.93 + -0.51 = -1.44
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"00111111111011100001010001111011"), -- 0.89 + 0.97 = 1.86
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"00111111110011100001010001111011"), -- 0.67 + 0.94 = 1.61
	(b"10111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111011001100110011001100110"), -- -0.32 + -0.58 = -0.9
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"10111111110010111000010100011110"), -- -0.77 + -0.82 = -1.59
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110101111010111000010100100", b"10111111100001010001111010111000"), -- -0.67 + -0.37 = -1.04
	(b"10111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111011010111000010100011111", b"10111111110000000000000000000000"), -- -0.58 + -0.92 = -1.5
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111101100110011001100110100"), -- 0.67 + 0.73 = 1.4
	(b"10111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110101011100001010001111011", b"10111111100000101000111101011100"), -- -0.68 + -0.34 = -1.02
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111111100000101000111101011100"), -- 0.23 + 0.79 = 1.02
	(b"10111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111011000010100011110101110", b"10111111101110011001100110011010"), -- -0.57 + -0.88 = -1.45
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111001101011100001010001111", b"10111111010000101000111101011100"), -- -0.05 + -0.71 = -0.76
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111011011100001010001111100"), -- -0.6 + -0.33 = -0.93
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111100001111010111000010100"), -- 0.17 + 0.89 = 1.06
	(b"00111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111111000000000000000000000000"), -- 0.45 + 0.05 = 0.5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111101111101011100001010010"), -- -0.7 + -0.79 = -1.49
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111101110000101000111101100"), -- 0.79 + 0.65 = 1.44
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"10111111010010100011110101110000"), -- -0.71 + -0.08 = -0.79
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111111101010111000010100011111"), -- 0.72 + 0.62 = 1.34
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111111000111000010100011110110"), -- 0.23 + 0.38 = 0.61
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111101111101011100001010001111", b"00111110100101000111101011100001"), -- 0.17 + 0.12 = 0.29
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111110110100011110101110000101"), -- -0.39 + -0.02 = -0.41
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111110110101110000101000111110"), -- -0.09 + -0.33 = -0.42
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"10111111100000010100011110101110"), -- -0.83 + -0.18 = -1.01
	(b"00111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"00111110111100001010001111010111"), -- 0.18 + 0.29 = 0.47
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111010111000010100011110110"), -- 0.62 + 0.24 = 0.86
	(b"10111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111101111000010100011110101110", b"10111111000001010001111010111000"), -- -0.41 + -0.11 = -0.52
	(b"10111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"10111111011110101110000101001000"), -- -0.94 + -0.04 = -0.98
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111110100011110101110000101001", b"10111111100100110011001100110011"), -- -0.87 + -0.28 = -1.15
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100101000111101011100001", b"10111110111000010100011110101110"), -- -0.15 + -0.29 = -0.44
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"00111111001000111101011100001010"), -- 0.36 + 0.28 = 0.64
	(b"00111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111000101000111101011100001"), -- 0.12 + 0.46 = 0.58
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000010100011110101110001", b"10111111101000000000000000000000"), -- -0.71 + -0.54 = -1.25
	(b"10111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111010101000111101011100001"), -- -0.21 + -0.62 = -0.83
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111001010001111010111000011", b"10111111101010100011110101110001"), -- -0.67 + -0.66 = -1.33
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"00111111011111010111000010100100"), -- 0 + 0.99 = 0.99
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111100001000111101011100001010", b"00111110101100110011001100110011"), -- 0.34 + 0.01 = 0.35
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"00111111010101110000101000111110"), -- 0.37 + 0.47 = 0.84
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111101100001010001111010111"), -- -0.76 + -0.62 = -1.38
	(b"10111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111010011001100110011001100"), -- -0.29 + -0.51 = -0.8
	(b"00111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111110010101110000101000111101"), -- 0.08 + 0.13 = 0.21
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111010111101011100001010010"), -- -0.67 + -0.2 = -0.87
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"00111111011000010100011110101110"), -- 0.43 + 0.45 = 0.88
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111011011100001010001111011"), -- -0.5 + -0.43 = -0.93
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"10111110001011100001010001111011"), -- -0.05 + -0.12 = -0.17
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111001010111000010100011110"), -- -0.26 + -0.41 = -0.67
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111001110000101000111101100", b"10111111100100110011001100110100"), -- -0.43 + -0.72 = -1.15
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111111101010100011110101110001"), -- 0.54 + 0.79 = 1.33
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"00111111100111000010100011110110"), -- 0.67 + 0.55 = 1.22
	(b"00111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111001010001111010111000011", b"00111111011100001010001111011000"), -- 0.28 + 0.66 = 0.94
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"10111111010000000000000000000000"), -- -0 + -0.75 = -0.75
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111010011110101110000101001"), -- -0.5 + -0.31 = -0.81
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110101011100001010001111011", b"10111111001100110011001100110100"), -- -0.36 + -0.34 = -0.7
	(b"10111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111100001010001111010111000"), -- -0.44 + -0.6 = -1.04
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111100100011110101110000110"), -- 0.54 + 0.6 = 1.14
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111010101110000101000111110"), -- 0.24 + 0.6 = 0.84
	(b"00111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111011110000101000111101100"), -- 0.09 + 0.88 = 0.97
	(b"00111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111111100011100001010001111011"), -- 0.68 + 0.43 = 1.11
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111101011100001010001111011"), -- -0.42 + -0.94 = -1.36
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111000010100011110101110001", b"10111111101011110101110000101001"), -- -0.83 + -0.54 = -1.37
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111011111010111000010100100"), -- -0.2 + -0.79 = -0.99
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111011110101110000101001000"), -- -0.65 + -0.33 = -0.98
	(b"00111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111111010100011110101110000101"), -- 0.68 + 0.14 = 0.82
	(b"00111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110110101110000101000111101", b"00111111101010100011110101110001"), -- 0.91 + 0.42 = 1.33
	(b"10111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111101110011001100110011010"), -- -0.55 + -0.9 = -1.45
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111000011110101110000101001", b"10111111101000000000000000000000"), -- -0.69 + -0.56 = -1.25
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111111000000000000000000000"), -- -0.96 + -0.79 = -1.75
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110101100110011001100110011", b"10111111011000010100011110101110"), -- -0.53 + -0.35 = -0.88
	(b"00111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111100010001111010111000010"), -- 0.53 + 0.54 = 1.07
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111011100110011001100110011", b"00111111110101011100001010010000"), -- 0.72 + 0.95 = 1.67
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"10111110101010001111010111000010"), -- -0.25 + -0.08 = -0.33
	(b"00111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111100001000111101011100001010", b"00111110110011001100110011001100"), -- 0.39 + 0.01 = 0.4
	(b"10111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111100111101011100001010010"), -- -0.29 + -0.95 = -1.24
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"10111111000000101000111101011100"), -- -0.04 + -0.47 = -0.51
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110110001111010111000010100", b"10111111100100110011001100110011"), -- -0.76 + -0.39 = -1.15
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"00111111101001010001111010111000"), -- 0.81 + 0.48 = 1.29
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111011100110011001100110011"), -- 0.3 + 0.65 = 0.95
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000101110000101000111101", b"00111111100110000101000111101100"), -- 0.6 + 0.59 = 1.19
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111011011100001010001111011", b"00111111101011100001010001111011"), -- 0.43 + 0.93 = 1.36
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110101000111101011100001010", b"10111110110100011110101110000101"), -- -0.09 + -0.32 = -0.41
	(b"10111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111011110000101000111101100"), -- -0.97 + -0 = -0.97
	(b"00111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110111010111000010100011110"), -- 0.26 + 0.2 = 0.46
	(b"10111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110110001111010111000010100", b"10111111001010001111010111000010"), -- -0.27 + -0.39 = -0.66
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111110000101000111101011100"), -- 0.79 + 0.73 = 1.52
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111011110101110000101001000", b"00111111101000000000000000000000"), -- 0.27 + 0.98 = 1.25
	(b"10111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111111011001100110011001100"), -- -0.95 + -0.9 = -1.85
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"00111111100011110101110000101001"), -- 0.25 + 0.87 = 1.12
	(b"00111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111000101110000101000111101", b"00111111010001010001111010111000"), -- 0.18 + 0.59 = 0.77
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"10111111000110011001100110011010"), -- -0.13 + -0.47 = -0.6
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111000001010001111010111000", b"10111111001100001010001111010111"), -- -0.17 + -0.52 = -0.69
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111011011100001010001111011", b"00111111100100110011001100110011"), -- 0.22 + 0.93 = 1.15
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111110111000010100011110110"), -- -0.77 + -0.95 = -1.72
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"10111110110000101000111101011100"), -- -0.16 + -0.22 = -0.38
	(b"00111110100111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111001011100001010001111011", b"00111111011111010111000010100100"), -- 0.31 + 0.68 = 0.99
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111100110000101000111101100"), -- -0.5 + -0.69 = -1.19
	(b"10111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111001101011100001010010000"), -- -0.38 + -0.33 = -0.71
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111001010001111010111000011", b"10111111101000101000111101011100"), -- -0.61 + -0.66 = -1.27
	(b"10111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111111010001111010111000010"), -- -0.98 + -0.84 = -1.82
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111100111101011100001010010"), -- -0.61 + -0.63 = -1.24
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"00111111101000010100011110101110"), -- 0.89 + 0.37 = 1.26
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111111100010001111010111000010"), -- 0.69 + 0.38 = 1.07
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"00111111100100110011001100110100"), -- 0.6 + 0.55 = 1.15
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"10111111010111101011100001010010"), -- -0.82 + -0.05 = -0.87
	(b"00111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111110010100011110101110000"), -- 0.75 + 0.83 = 1.58
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"10111111100010111000010100011111"), -- -0.87 + -0.22 = -1.09
	(b"00111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111001100001010001111010111", b"00111111110000101000111101011100"), -- 0.83 + 0.69 = 1.52
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111000111000010100011110110", b"00111111100111010111000010100100"), -- 0.62 + 0.61 = 1.23
	(b"10111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111100101000111101011100001"), -- -0.46 + -0.7 = -1.16
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"10111110100001010001111010111000"), -- -0.09 + -0.17 = -0.26
	(b"10111110100111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"10111110111110101110000101001000"), -- -0.31 + -0.18 = -0.49
	(b"10111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111100110011001100110011010"), -- -0.56 + -0.64 = -1.2
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"00111111011001100110011001100110"), -- 0.35 + 0.55 = 0.9
	(b"10111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111001010111000010100011111", b"10111111100000000000000000000000"), -- -0.33 + -0.67 = -1
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111110101011100001010001111011"), -- -0.15 + -0.19 = -0.34
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111110101000111101011100001010", b"10111111001100001010001111010111"), -- -0.37 + -0.32 = -0.69
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111100100001010001111010111"), -- -0.26 + -0.87 = -1.13
	(b"00111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111100000010100011110101110"), -- 0.61 + 0.4 = 1.01
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"10111111000110011001100110011010"), -- -0.54 + -0.06 = -0.6
	(b"10111111011011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111111101001111010111000010100"), -- -0.93 + -0.38 = -1.31
	(b"10111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111001011100001010001111011", b"10111111110100110011001100110100"), -- -0.97 + -0.68 = -1.65
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111101101110000101000111101100", b"10111111011001100110011001100110"), -- -0.81 + -0.09 = -0.9
	(b"00111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111001111010111000010100100", b"00111111100101000111101011100001"), -- 0.42 + 0.74 = 1.16
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111001110000101000111101100", b"00111111011100001010001111011000"), -- 0.22 + 0.72 = 0.94
	(b"00111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111100011100001010001111011"), -- 0.65 + 0.46 = 1.11
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"00111111101100001010001111010111"), -- 0.54 + 0.84 = 1.38
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"10111111100001111010111000010100"), -- -0.89 + -0.17 = -1.06
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111101011100001010001111011"), -- 0.55 + 0.81 = 1.36
	(b"10111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111110101011100001010001111011", b"10111111010000000000000000000000"), -- -0.41 + -0.34 = -0.75
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111101001111010111000010100"), -- -0.67 + -0.64 = -1.31
	(b"10111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"10111111101011001100110011001101"), -- -0.91 + -0.44 = -1.35
	(b"00111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111000110011001100110011010"), -- 0.06 + 0.54 = 0.6
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110100010100011110101110001", b"10111111100111010111000010100100"), -- -0.96 + -0.27 = -1.23
	(b"00111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110101110000101000111101100", b"00111111011110000101000111101100"), -- 0.61 + 0.36 = 0.97
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111100110101110000101001000"), -- -0.8 + -0.41 = -1.21
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"10111111101100110011001100110100"), -- -0.49 + -0.91 = -1.4
	(b"00111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111111000000000000000000000"), -- 0.85 + 0.9 = 1.75
	(b"00111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"00111111000101000111101011100001"), -- 0.19 + 0.39 = 0.58
	(b"00111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111000011110101110000101001", b"00111111101100001010001111010111"), -- 0.82 + 0.56 = 1.38
	(b"00111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111001001100110011001100110"), -- 0.07 + 0.58 = 0.65
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111010001010001111010111000", b"10111111101111010111000010100100"), -- -0.71 + -0.77 = -1.48
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111100000000000000000000000"), -- 0.8 + 0.2 = 1
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111101011001100110011001100"), -- 0.52 + 0.83 = 1.35
	(b"00111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110111000010100011110101110", b"00111111000100011110101110000101"), -- 0.13 + 0.44 = 0.57
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111100011001100110011001101"), -- -0.79 + -0.31 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"00111101011101011100001010001111"), -- 0 + 0.06 = 0.06
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"00111111100001010001111010111000"), -- 0.59 + 0.45 = 1.04
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111101111000010100011110110"), -- -0.84 + -0.63 = -1.47
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"00111111110001111010111000010100"), -- 0.72 + 0.84 = 1.56
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111011010001111010111000011", b"00111111100101110000101000111110"), -- 0.27 + 0.91 = 1.18
	(b"10111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111111010110011001100110011010"), -- -0.66 + -0.19 = -0.85
	(b"00111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111100110011001100110011010"), -- 0.39 + 0.81 = 1.2
	(b"10111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111010011110101110000101001", b"10111111100000000000000000000000"), -- -0.19 + -0.81 = -1
	(b"00111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"00111110011010111000010100011111"), -- 0.06 + 0.17 = 0.23
	(b"10111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111000111101011100001010010"), -- -0.29 + -0.33 = -0.62
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111001010111000010100011111"), -- -0.04 + -0.63 = -0.67
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111111101000000000000000000000"), -- -0.8 + -0.45 = -1.25
	(b"00111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"00111111011101011100001010010000"), -- 0.92 + 0.04 = 0.96
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111111001100001010001111010111"), -- 0.56 + 0.13 = 0.69
	(b"10111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111100100011110101110000101"), -- -0.56 + -0.58 = -1.14
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111011110101110000101001000", b"00111111101101000111101011100010"), -- 0.43 + 0.98 = 1.41
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010000101000111101011100", b"10111111101110101110000101001000"), -- -0.7 + -0.76 = -1.46
	(b"00111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111000001111010111000010100", b"00111111100001111010111000010100"), -- 0.53 + 0.53 = 1.06
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111101110011001100110011010"), -- 0.95 + 0.5 = 1.45
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"10111111100001111010111000010100"), -- -0.23 + -0.83 = -1.06
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111101010100011110101110000"), -- -0.69 + -0.64 = -1.33
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111101001010001111010111000"), -- -0.65 + -0.64 = -1.29
	(b"10111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"10111111000110011001100110011010"), -- -0.34 + -0.26 = -0.6
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111101001010001111010111000"), -- 0.79 + 0.5 = 1.29
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111101011001100110011001100"), -- -0.76 + -0.59 = -1.35
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"00111111011110101110000101001000"), -- 0.5 + 0.48 = 0.98
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011110101110000101001000", b"10111111011110101110000101001000"), -- -0 + -0.98 = -0.98
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111010000101000111101011100"), -- 0.27 + 0.49 = 0.76
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"10111111011001100110011001100110"), -- -0.43 + -0.47 = -0.9
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"00111111001100001010001111010111"), -- 0.52 + 0.17 = 0.69
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011101011100001010001111", b"00111111100101000111101011100001"), -- 0.2 + 0.96 = 1.16
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111001100110011001100110011"), -- -0.39 + -0.31 = -0.7
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111100110011001100110011010"), -- -0.8 + -0.4 = -1.2
	(b"10111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111100000010100011110101110"), -- -0.58 + -0.43 = -1.01
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111010001111010111000010100"), -- -0.48 + -0.3 = -0.78
	(b"00111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111010000101000111101011100"), -- 0.03 + 0.73 = 0.76
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111011100110011001100110011", b"00111111100011110101110000101001"), -- 0.17 + 0.95 = 1.12
	(b"00111110111100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111111000001010001111010111000"), -- 0.47 + 0.05 = 0.52
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001110101110000101001000", b"10111111110110000101000111101100"), -- -0.96 + -0.73 = -1.69
	(b"00111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111101111000010100011110101110", b"00111111000001111010111000010100"), -- 0.42 + 0.11 = 0.53
	(b"10111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111100001111010111000010100"), -- -0.63 + -0.43 = -1.06
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111010000000000000000000000", b"00111111101111000010100011110110"), -- 0.72 + 0.75 = 1.47
	(b"00111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111100101000111101011100001010", b"00111110111010111000010100011111"), -- 0.44 + 0.02 = 0.46
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111111100001100110011001100110"), -- 0.89 + 0.16 = 1.05
	(b"10111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"10111110100110011001100110011010"), -- -0.08 + -0.22 = -0.3
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110000001010001111010111000", b"10111111001001100110011001100110"), -- -0.52 + -0.13 = -0.65
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"10111111100000101000111101011100"), -- -0.96 + -0.06 = -1.02
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"00111111000111101011100001010010"), -- 0.43 + 0.19 = 0.62
	(b"10111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111101111000010100011110101110", b"10111110100101000111101011100010"), -- -0.18 + -0.11 = -0.29
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110110101110000101000111101", b"10111111001011100001010001111010"), -- -0.26 + -0.42 = -0.68
	(b"00111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"00111110111010111000010100011111"), -- 0.09 + 0.37 = 0.46
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110110101110000101000111101", b"10111111001010001111010111000010"), -- -0.24 + -0.42 = -0.66
	(b"10111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111111101110000101000111110"), -- -0.94 + -0.99 = -1.93
	(b"10111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"10111111100001111010111000010101"), -- -0.21 + -0.85 = -1.06
	(b"10111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"10111111100000010100011110101110"), -- -0.95 + -0.06 = -1.01
	(b"00111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111000100011110101110000101", b"00111111011110101110000101001000"), -- 0.41 + 0.57 = 0.98
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"10111110101011100001010001111011"), -- -0.3 + -0.04 = -0.34
	(b"00111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111011000111101011100001010"), -- 0.08 + 0.81 = 0.89
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110000001010001111010111000", b"10111110110100011110101110000101"), -- -0.28 + -0.13 = -0.41
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111100101011100001010001111"), -- -0.64 + -0.53 = -1.17
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111110111110101110000101001000"), -- 0.36 + 0.13 = 0.49
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111111100000101000111101011100"), -- 0.23 + 0.79 = 1.02
	(b"00111111011011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"00111111101100110011001100110011"), -- 0.93 + 0.47 = 1.4
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111110100011110101110000101"), -- 0.81 + 0.83 = 1.64
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111110010001111010111000010"), -- 0.69 + 0.88 = 1.57
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111010001010001111010111000"), -- 0.25 + 0.52 = 0.77
	(b"10111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"10111111111100011110101110000110"), -- -0.98 + -0.91 = -1.89
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111100000101000111101011100"), -- -0.39 + -0.63 = -1.02
	(b"00111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111101100001010001111010111"), -- 0.48 + 0.9 = 1.38
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"00111111001100001010001111010111"), -- 0.22 + 0.47 = 0.69
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111010011110101110000101001"), -- -0.24 + -0.57 = -0.81
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111100110011001100110011010"), -- 0.74 + 0.46 = 1.2
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"00111111001011100001010001111011"), -- 0.62 + 0.06 = 0.68
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111100101011100001010001111"), -- -0.53 + -0.64 = -1.17
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"10111110010101110000101000111110"), -- -0.17 + -0.04 = -0.21
	(b"00111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011011100001010001111011", b"00111111100001100110011001100110"), -- 0.12 + 0.93 = 1.05
	(b"00111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111000111000010100011110110", b"00111111101110011001100110011010"), -- 0.84 + 0.61 = 1.45
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111011011100001010001111011"), -- 0.05 + 0.88 = 0.93
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010001010001111010111000", b"10111111100010001111010111000010"), -- -0.3 + -0.77 = -1.07
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111100111010111000010100100"), -- 0.74 + 0.49 = 1.23
	(b"00111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111001110000101000111101100", b"00111111011110101110000101001000"), -- 0.26 + 0.72 = 0.98
	(b"10111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111100010100011110101110001"), -- -0.21 + -0.87 = -1.08
	(b"10111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"10111111000101000111101011100001"), -- -0.11 + -0.47 = -0.58
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111010100011110101110000101", b"00111111101100011110101110000101"), -- 0.57 + 0.82 = 1.39
	(b"00111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"00111110110100011110101110000101"), -- 0.19 + 0.22 = 0.41
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010000101000111101011100", b"10111111101101110000101000111110"), -- -0.67 + -0.76 = -1.43
	(b"00111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"00111111000011001100110011001101"), -- 0.07 + 0.48 = 0.55
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111110011110101110000101001"), -- -0.82 + -0.8 = -1.62
	(b"10111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111100000000000000000000000"), -- -0.41 + -0.59 = -1
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101111000010100011110101110", b"10111111000011110101110000101001"), -- -0.45 + -0.11 = -0.56
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111100111101011100001010010"), -- 0.57 + 0.67 = 1.24
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111010110011001100110011010"), -- -0.28 + -0.57 = -0.85
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110111010111000010100011111", b"10111111011111010111000010100100"), -- -0.53 + -0.46 = -0.99
	(b"10111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001110101110000101001000", b"10111111100010100011110101110001"), -- -0.35 + -0.73 = -1.08
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"10111111100000000000000000000000"), -- -0.25 + -0.75 = -1
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"10111111100000010100011110101110"), -- -0.26 + -0.75 = -1.01
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111111000011001100110011001101"), -- -0.1 + -0.45 = -0.55
	(b"10111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111110100010100011110101110001", b"10111111100000000000000000000000"), -- -0.73 + -0.27 = -1
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111011101011100001010001111"), -- -0.37 + -0.59 = -0.96
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"00111111000000101000111101011100"), -- 0.22 + 0.29 = 0.51
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111100011001100110011001101"), -- 0.5 + 0.6 = 1.1
	(b"10111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111100000010100011110101110"), -- -0.02 + -0.99 = -1.01
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111010011001100110011001101"), -- 0.2 + 0.6 = 0.8
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"10111111101111101011100001010010"), -- -0.6 + -0.89 = -1.49
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111100101011100001010001111"), -- 0.52 + 0.65 = 1.17
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"10111111011100001010001111010111"), -- -0.8 + -0.14 = -0.94
	(b"10111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"10111111101011110101110000101001"), -- -0.63 + -0.74 = -1.37
	(b"00111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"00111111011110000101000111101100"), -- 0.66 + 0.31 = 0.97
	(b"00111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111010111000010100011110110", b"00111111111000101000111101011100"), -- 0.91 + 0.86 = 1.77
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"10111110001000111101011100001010"), -- -0.1 + -0.06 = -0.16
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111010000000000000000000000"), -- -0.17 + -0.58 = -0.75
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111010011001100110011001100"), -- 0.22 + 0.58 = 0.8
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111101000010100011110101110"), -- 0.74 + 0.52 = 1.26
	(b"10111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"10111111010001111010111000010101"), -- -0.73 + -0.05 = -0.78
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001011100001010001111011", b"10111111011011100001010001111011"), -- -0.25 + -0.68 = -0.93
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001110000101000111101100", b"00111111100000101000111101011100"), -- 0.3 + 0.72 = 1.02
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"10111111101111000010100011110110"), -- -0.69 + -0.78 = -1.47
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111010110011001100110011010", b"00111111110010100011110101110001"), -- 0.73 + 0.85 = 1.58
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111001000010100011110101110", b"00111111101110000101000111101100"), -- 0.81 + 0.63 = 1.44
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111111001110101110000101000111"), -- 0.59 + 0.14 = 0.73
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111100111000010100011110110"), -- 0.73 + 0.49 = 1.22
	(b"10111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110100000000000000000000000", b"10111111011000010100011110101110"), -- -0.63 + -0.25 = -0.88
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111110010111000010100011111"), -- 0.86 + 0.73 = 1.59
	(b"00111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111111100000101000111101011100"), -- 0.94 + 0.08 = 1.02
	(b"10111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"10111111111010111000010100011110"), -- -0.88 + -0.96 = -1.84
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111110101011100001010010000"), -- 0.86 + 0.81 = 1.67
	(b"00111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"00111111011101011100001010010000"), -- 0.41 + 0.55 = 0.96
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111101011100001010001111011"), -- 0.56 + 0.8 = 1.36
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111100101000111101011100001"), -- -0.76 + -0.4 = -1.16
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111101100011110101110000101001"), -- -0.05 + -0.02 = -0.07
	(b"00111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111111101110101110000101001000"), -- 0.84 + 0.62 = 1.46
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"00111110110000101000111101011100"), -- 0.34 + 0.04 = 0.38
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111111100000101000111101011100"), -- 0.59 + 0.43 = 1.02
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011010111000010100011111", b"00111111011011100001010001111011"), -- 0.01 + 0.92 = 0.93
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111111100001111010111000010100"), -- 0.63 + 0.43 = 1.06
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111011010111000010100011111"), -- 0.43 + 0.49 = 0.92
	(b"10111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"10111110100010100011110101110001"), -- -0.22 + -0.05 = -0.27
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110101011100001010001111011", b"10111110110011001100110011001101"), -- -0.06 + -0.34 = -0.4
	(b"00111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111000110011001100110011001"), -- 0.08 + 0.52 = 0.6
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111100101110000101000111110"), -- -0.67 + -0.51 = -1.18
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111101001010001111010111000"), -- -0.49 + -0.8 = -1.29
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111001111010111000010100100", b"00111111110110101110000101001000"), -- 0.97 + 0.74 = 1.71
	(b"00111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111111010001111010111000010100"), -- 0.64 + 0.14 = 0.78
	(b"00111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011110101110000101001000", b"00111111111110000101000111101100"), -- 0.96 + 0.98 = 1.94
	(b"10111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"10111111010001111010111000010101"), -- -0.66 + -0.12 = -0.78
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"10111111100101011100001010010000"), -- -0.26 + -0.91 = -1.17
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111000000101000111101011100", b"00111111001110000101000111101011"), -- 0.21 + 0.51 = 0.72
	(b"10111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111100111000010100011110110"), -- -0.62 + -0.6 = -1.22
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010110011001100110011010", b"00111111100010100011110101110001"), -- 0.23 + 0.85 = 1.08
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"00111110111110101110000101001000"), -- 0.2 + 0.29 = 0.49
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111100011100001010001111011"), -- -0.6 + -0.51 = -1.11
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"10111111101010001111010111000010"), -- -0.5 + -0.82 = -1.32
	(b"10111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111000000101000111101011100"), -- -0.18 + -0.33 = -0.51
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111010001111010111000010100"), -- 0.38 + 0.4 = 0.78
	(b"00111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111111011110000101000111101100"), -- 0.18 + 0.79 = 0.97
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110110101110000101000111101", b"00111111010011001100110011001100"), -- 0.38 + 0.42 = 0.8
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111000010100011110101110001"), -- -0.54 + -0 = -0.54
	(b"00111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"00111111100010001111010111000010"), -- 0.88 + 0.19 = 1.07
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111001101011100001010010000"), -- 0.25 + 0.46 = 0.71
	(b"10111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111111101100110011001100110011"), -- -0.95 + -0.45 = -1.4
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111100000010100011110101110"), -- 0.52 + 0.49 = 1.01
	(b"10111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111111000111101011100001010"), -- -0.91 + -0.87 = -1.78
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111101010100011110101110000"), -- -0.83 + -0.5 = -1.33
	(b"00111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111010001111010111000010101"), -- 0.11 + 0.67 = 0.78
	(b"10111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111100010111000010100011111"), -- -0.68 + -0.41 = -1.09
	(b"10111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110000001010001111010111000", b"10111110100000000000000000000000"), -- -0.12 + -0.13 = -0.25
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111110110100011110101110000101"), -- 0.25 + 0.16 = 0.41
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111011110101110000101001000"), -- 0.34 + 0.64 = 0.98
	(b"00111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"00111111101110101110000101001000"), -- 0.99 + 0.47 = 1.46
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111100011110101110000101001"), -- -0.81 + -0.31 = -1.12
	(b"10111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"10111111001100001010001111010111"), -- -0.66 + -0.03 = -0.69
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111100001000111101011100001010", b"00111110110001111010111000010100"), -- 0.38 + 0.01 = 0.39
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111000100011110101110000101"), -- 0.17 + 0.4 = 0.57
	(b"00111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111011101011100001010001111", b"00111111111011110101110000101001"), -- 0.91 + 0.96 = 1.87
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111100001100110011001100110"), -- 0.38 + 0.67 = 1.05
	(b"00111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111001000010100011110101110", b"00111111101110101110000101001000"), -- 0.83 + 0.63 = 1.46
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111010000101000111101011100", b"10111111101110011001100110011010"), -- -0.69 + -0.76 = -1.45
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111010001010001111010111000", b"10111111010111000010100011110110"), -- -0.09 + -0.77 = -0.86
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110101100110011001100110011", b"10111111001111010111000010100100"), -- -0.39 + -0.35 = -0.74
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110110101110000101000111101", b"10111111010001111010111000010100"), -- -0.36 + -0.42 = -0.78
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111010010100011110101110001"), -- -0.36 + -0.43 = -0.79
	(b"00111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"00111111111011100001010001111011"), -- 0.92 + 0.94 = 1.86
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"10111110011000010100011110101110"), -- -0.06 + -0.16 = -0.22
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111110010111000010100011110"), -- -0.65 + -0.94 = -1.59
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111101110000101000111101100"), -- -0.82 + -0.62 = -1.44
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001111010111000010100100"), -- 0.04 + 0.7 = 0.74
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000111000010100011110110", b"00111111100011100001010001111011"), -- 0.5 + 0.61 = 1.11
	(b"00111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000011110101110000101001", b"00111111100110101110000101001000"), -- 0.65 + 0.56 = 1.21
	(b"00111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111111100010100011110101110000"), -- 0.65 + 0.43 = 1.08
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111010100011110101110000110"), -- -0.72 + -0.1 = -0.82
	(b"00111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111010100011110101110000101", b"00111111100000000000000000000000"), -- 0.18 + 0.82 = 1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"10111111011000010100011110101110"), -- -0.7 + -0.18 = -0.88
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110011010111000010100011111", b"10111111000001111010111000010101"), -- -0.3 + -0.23 = -0.53
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111100011001100110011001100"), -- -0.26 + -0.84 = -1.1
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111101101110000101000111101100", b"10111110000001010001111010111000"), -- -0.04 + -0.09 = -0.13
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111010100011110101110000101"), -- 0.17 + 0.65 = 0.82
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111111000000000000000000000000"), -- 0.37 + 0.13 = 0.5
	(b"10111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"10111111010001010001111010111000"), -- -0.51 + -0.26 = -0.77
	(b"00111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"00111111010011110101110000101001"), -- 0.48 + 0.33 = 0.81
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"10111111001111010111000010100100"), -- -0.52 + -0.22 = -0.74
	(b"00111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111010000000000000000000000"), -- 0.45 + 0.3 = 0.75
	(b"00111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111011000111101011100001010"), -- 0.39 + 0.5 = 0.89
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"10111111100000010100011110101110"), -- -0.89 + -0.12 = -1.01
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111010011001100110011001101"), -- 0.56 + 0.24 = 0.8
	(b"10111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111101110101110000101001000"), -- -0.95 + -0.51 = -1.46
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111101001100110011001100110"), -- 0.9 + 0.4 = 1.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110111101011100001010001111", b"10111111001011100001010001111011"), -- -0.2 + -0.48 = -0.68
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"10111111110010100011110101110000"), -- -0.8 + -0.78 = -1.58
	(b"10111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111110101111010111000010100100", b"10111111101011001100110011001101"), -- -0.98 + -0.37 = -1.35
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111100100110011001100110011"), -- 0.35 + 0.8 = 1.15
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111100111000010100011110110"), -- -0.64 + -0.58 = -1.22
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"10111111011101011100001010001111"), -- -0.82 + -0.14 = -0.96
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111110100110011001100110011"), -- -0.81 + -0.84 = -1.65
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"00111110011010111000010100011111"), -- 0.01 + 0.22 = 0.23
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"00111101101000111101011100001010"), -- 0.04 + 0.04 = 0.08
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111100001010001111010111000"), -- -0.45 + -0.59 = -1.04
	(b"00111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111011110101110000101001000"), -- 0.15 + 0.83 = 0.98
	(b"00111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111101010001111010111000011"), -- 0.92 + 0.4 = 1.32
	(b"00111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"00111111110011001100110011001101"), -- 0.66 + 0.94 = 1.6
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111101111000010100011110101110", b"10111111010111101011100001010010"), -- -0.76 + -0.11 = -0.87
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"10111110110111000010100011110101"), -- -0.39 + -0.04 = -0.43
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110111110101110000101001000", b"10111111100110011001100110011010"), -- -0.71 + -0.49 = -1.2
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110101100110011001100110011", b"10111111101001111010111000010100"), -- -0.96 + -0.35 = -1.31
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"10111111101000101000111101011100"), -- -0.36 + -0.91 = -1.27
	(b"10111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111000101110000101000111101"), -- -0.08 + -0.51 = -0.59
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111001100001010001111010111", b"00111111010111000010100011110110"), -- 0.17 + 0.69 = 0.86
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"00111111001101011100001010010000"), -- 0.43 + 0.28 = 0.71
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"00111111101001111010111000010100"), -- 0.32 + 0.99 = 1.31
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"00111110110101110000101000111101"), -- 0.35 + 0.07 = 0.42
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111000111101011100001010010"), -- 0.22 + 0.4 = 0.62
	(b"00111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011100110011001100110011", b"00111111100011001100110011001101"), -- 0.15 + 0.95 = 1.1
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111111100011110101110000101001"), -- 0.5 + 0.62 = 1.12
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111001101011100001010010000"), -- -0.09 + -0.62 = -0.71
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111011011100001010001111011", b"10111111101110101110000101001000"), -- -0.53 + -0.93 = -1.46
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"00111111001110101110000101000111"), -- 0.7 + 0.03 = 0.73
	(b"00111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"00111111010001111010111000010101"), -- 0.61 + 0.17 = 0.78
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110111110101110000101001000", b"10111111000010100011110101110001"), -- -0.05 + -0.49 = -0.54
	(b"00111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"00111111101110000101000111101100"), -- 0.99 + 0.45 = 1.44
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"00111111000101110000101000111110"), -- 0.3 + 0.29 = 0.59
	(b"10111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"10111110011000010100011110101110"), -- -0.08 + -0.14 = -0.22
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110111100001010001111011000"), -- 0.17 + 0.3 = 0.47
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111101000000000000000000000"), -- -0.67 + -0.58 = -1.25
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111000010100011110101110001", b"10111111101101000111101011100010"), -- -0.87 + -0.54 = -1.41
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111100111010111000010100100"), -- 0.4 + 0.83 = 1.23
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110100101000111101011100001", b"10111111001110000101000111101100"), -- -0.43 + -0.29 = -0.72
	(b"00111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111101011001100110011001101"), -- 0.85 + 0.5 = 1.35
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111011110000101000111101100", b"10111111101111101011100001010010"), -- -0.52 + -0.97 = -1.49
	(b"10111110111100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111101110101110000101001000"), -- -0.47 + -0.99 = -1.46
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"10111111110011100001010001111011"), -- -0.86 + -0.75 = -1.61
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111111010110011001100110011001"), -- -0.83 + -0.02 = -0.85
	(b"00111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"00111111001010001111010111000011"), -- 0.33 + 0.33 = 0.66
	(b"00111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111001010001111010111000011", b"00111111100010100011110101110001"), -- 0.42 + 0.66 = 1.08
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111010111000010100011110110"), -- 0.34 + 0.52 = 0.86
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"00111101010011001100110011001100"), -- 0.02 + 0.03 = 0.05
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"00111110111101011100001010001111"), -- 0 + 0.48 = 0.48
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111101010100011110101110001"), -- -0.92 + -0.41 = -1.33
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"10111111001011100001010001111011"), -- -0.54 + -0.14 = -0.68
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111010110011001100110011010"), -- 0.36 + 0.49 = 0.85
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111001110000101000111101100", b"00111111011111010111000010100100"), -- 0.27 + 0.72 = 0.99
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111001110101110000101001000"), -- -0.15 + -0.58 = -0.73
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011000010100011110101110", b"10111111110010100011110101110000"), -- -0.7 + -0.88 = -1.58
	(b"00111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111000111101011100001010010"), -- 0.42 + 0.2 = 0.62
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111101001100110011001100110"), -- -0.72 + -0.58 = -1.3
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"10111111100000000000000000000000"), -- -0.84 + -0.16 = -1
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111011110101110000101000111"), -- -0.45 + -0.53 = -0.98
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"10111111101101000111101011100010"), -- -0.5 + -0.91 = -1.41
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111000011001100110011001101", b"10111111100010100011110101110000"), -- -0.53 + -0.55 = -1.08
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111100110011001100110011010"), -- -0.36 + -0.84 = -1.2
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111110001010001111010111000"), -- 0.74 + 0.8 = 1.54
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110011010111000010100011111", b"10111111011000010100011110101110"), -- -0.65 + -0.23 = -0.88
	(b"10111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111111000111101011100001010"), -- -0.99 + -0.79 = -1.78
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111101100001010001111010111"), -- -0.76 + -0.62 = -1.38
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111111100001100110011001100110"), -- -0.86 + -0.19 = -1.05
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111111010000000000000000000000"), -- 0.37 + 0.38 = 0.75
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"10111111100000000000000000000000"), -- -0.86 + -0.14 = -1
	(b"10111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111110101110000101000111110"), -- -0.88 + -0.8 = -1.68
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110110101110000101000111101", b"10111111100110000101000111101011"), -- -0.77 + -0.42 = -1.19
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111011101011100001010001111"), -- 0.32 + 0.64 = 0.96
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111111000100011110101110000101"), -- 0.57 + 0 = 0.57
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111011110000101000111101100"), -- -0.64 + -0.33 = -0.97
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001011100001010001111011", b"10111111001111010111000010100100"), -- -0.06 + -0.68 = -0.74
	(b"00111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"00111110110001111010111000010101"), -- 0.06 + 0.33 = 0.39
	(b"10111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111101011100001010001111011"), -- -0.57 + -0.79 = -1.36
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111011100110011001100110100"), -- 0.35 + 0.6 = 0.95
	(b"00111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111110010001111010111000010"), -- 0.68 + 0.89 = 1.57
	(b"00111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111101001111010111000010100"), -- 0.42 + 0.89 = 1.31
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111000011001100110011001101"), -- 0.25 + 0.3 = 0.55
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111111001100001010001111010111"), -- 0.69 + 0 = 0.69
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111011101011100001010010000"), -- 0.23 + 0.73 = 0.96
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"00111111100011100001010001111011"), -- 0.72 + 0.39 = 1.11
	(b"00111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111011111010111000010100100"), -- 0.49 + 0.5 = 0.99
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111010011001100110011001101"), -- -0.3 + -0.5 = -0.8
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111111010111101011100001010010"), -- -0.42 + -0.45 = -0.87
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111110101000111101011100001011"), -- -0.3 + -0.02 = -0.32
	(b"00111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111100101000111101011100001010", b"00111111010101110000101000111101"), -- 0.82 + 0.02 = 0.84
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"10111111000000000000000000000000"), -- -0.06 + -0.44 = -0.5
	(b"00111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111100101011100001010001111"), -- 0.77 + 0.4 = 1.17
	(b"10111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111011101011100001010010000"), -- -0.27 + -0.69 = -0.96
	(b"10111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110101100110011001100110011", b"10111111100011001100110011001101"), -- -0.75 + -0.35 = -1.1
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111000111101011100001010010"), -- -0.09 + -0.53 = -0.62
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"10111110111100001010001111010110"), -- -0.39 + -0.08 = -0.47
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"10111111101000000000000000000000"), -- -0.78 + -0.47 = -1.25
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111011011100001010001111011"), -- 0.05 + 0.88 = 0.93
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- -0 + -0.3 = -0.3
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111101111000010100011110101110", b"10111110111101011100001010010000"), -- -0.37 + -0.11 = -0.48
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010111000010100011110110", b"00111111010111000010100011110110"), -- 0 + 0.86 = 0.86
	(b"00111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"00111111100011110101110000101001"), -- 0.75 + 0.37 = 1.12
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"00111110110101110000101000111110"), -- 0.17 + 0.25 = 0.42
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"00111111100000111101011100001010"), -- 0.55 + 0.48 = 1.03
	(b"10111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111110100101000111101011100001", b"10111111100000111101011100001010"), -- -0.74 + -0.29 = -1.03
	(b"00111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"00111111111011100001010001111011"), -- 0.87 + 0.99 = 1.86
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"10111111111001100110011001100110"), -- -0.84 + -0.96 = -1.8
	(b"10111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111011001100110011001100110"), -- -0.03 + -0.87 = -0.9
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110110001111010111000010100", b"10111111010001111010111000010100"), -- -0.39 + -0.39 = -0.78
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"00111110100101000111101011100001"), -- 0.04 + 0.25 = 0.29
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111011100001010001111010111"), -- -0.84 + -0.1 = -0.94
	(b"10111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111111101011100001010010000"), -- -0.97 + -0.95 = -1.92
	(b"00111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"00111110111110101110000101000111"), -- 0.42 + 0.07 = 0.49
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111110111101011100001010010"), -- -0.8 + -0.94 = -1.74
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111101101110000101000111101100", b"00111111001101011100001010010000"), -- 0.62 + 0.09 = 0.71
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111110100001010001111010111000"), -- 0.1 + 0.16 = 0.26
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111000011110101110000101001", b"10111111001110101110000101001000"), -- -0.17 + -0.56 = -0.73
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110111010111000010100011111", b"10111111010100011110101110000110"), -- -0.36 + -0.46 = -0.82
	(b"00111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110001110000101000111101100", b"00111110100000000000000000000000"), -- 0.07 + 0.18 = 0.25
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"00111111110111010111000010100100"), -- 0.89 + 0.84 = 1.73
	(b"00111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111110011110101110000101001"), -- 0.98 + 0.64 = 1.62
	(b"00111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111000111101011100001010010"), -- 0.13 + 0.49 = 0.62
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111111010010100011110101110001"), -- 0.79 + 0 = 0.79
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111010000000000000000000000", b"00111111110000111101011100001010"), -- 0.78 + 0.75 = 1.53
	(b"10111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"10111110110111000010100011110110"), -- -0.29 + -0.14 = -0.43
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111001100110011001100110100"), -- -0.1 + -0.6 = -0.7
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111011000111101011100001011"), -- -0.1 + -0.79 = -0.89
	(b"00111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111100100110011001100110011"), -- 0.48 + 0.67 = 1.15
	(b"00111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111110010000101000111101011100"), -- 0.11 + 0.08 = 0.19
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111001010111000010100011111", b"10111111001011100001010001111011"), -- -0.01 + -0.67 = -0.68
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111011101011100001010010000"), -- 0.5 + 0.46 = 0.96
	(b"00111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110101110000101000111101100", b"00111111100010001111010111000010"), -- 0.71 + 0.36 = 1.07
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111100111101011100001010010"), -- -0.4 + -0.84 = -1.24
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111101110011001100110011010"), -- 0.78 + 0.67 = 1.45
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"00111111100101110000101000111101"), -- 0.24 + 0.94 = 1.18
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111100010100011110101110000"), -- 0.38 + 0.7 = 1.08
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110001110000101000111101100", b"00111111100100110011001100110100"), -- 0.97 + 0.18 = 1.15
	(b"00111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111111000111000010100011110110"), -- 0.61 + 0 = 0.61
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111111100001010001111010111"), -- -0.89 + -0.99 = -1.88
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"00111111100101000111101011100001"), -- 0.17 + 0.99 = 1.16
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"10111111011111010111000010100011"), -- -0.96 + -0.03 = -0.99
	(b"00111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111100000101000111101011100"), -- 0.44 + 0.58 = 1.02
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111100111010111000010100100"), -- 0.69 + 0.54 = 1.23
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111101011001100110011001101"), -- 0.95 + 0.4 = 1.35
	(b"00111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111110101011100001010001111"), -- 0.84 + 0.83 = 1.67
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111000101110000101000111101"), -- 0.35 + 0.24 = 0.59
	(b"10111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000011110101110000101001", b"10111111011010001111010111000010"), -- -0.35 + -0.56 = -0.91
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110111110101110000101001000", b"10111111001111010111000010100100"), -- -0.25 + -0.49 = -0.74
	(b"10111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111101100001010001111010111"), -- -0.44 + -0.94 = -1.38
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111111000010100011110101110"), -- -0.77 + -0.99 = -1.76
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"10111110001110000101000111101100"), -- -0.15 + -0.03 = -0.18
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111111101001100110011001100110"), -- -0.92 + -0.38 = -1.3
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111110000111101011100001010"), -- -0.96 + -0.57 = -1.53
	(b"10111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110100000000000000000000000", b"10111110101000111101011100001010"), -- -0.07 + -0.25 = -0.32
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"00111110100001010001111010111000"), -- 0.2 + 0.06 = 0.26
	(b"00111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110101110000101000111101100", b"00111111100001010001111010111000"), -- 0.68 + 0.36 = 1.04
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"10111111110010100011110101110000"), -- -0.69 + -0.89 = -1.58
	(b"00111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111111100011001100110011001101"), -- 0.48 + 0.62 = 1.1
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111111011010001111010111000010"), -- 0.29 + 0.62 = 0.91
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111111001110000101000111101100"), -- 0.29 + 0.43 = 0.72
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111011010111000010100011111", b"00111111111100011110101110000110"), -- 0.97 + 0.92 = 1.89
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111111001110000101000111101011"), -- -0.7 + -0.02 = -0.72
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111101001111010111000010101"), -- 0.97 + 0.34 = 1.31
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110101100110011001100110011", b"10111111100101000111101011100001"), -- -0.81 + -0.35 = -1.16
	(b"10111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111101100011110101110000101001"), -- -0.07 + -0 = -0.07
	(b"10111110100111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111110101111010111000010100100", b"10111111001011100001010001111011"), -- -0.31 + -0.37 = -0.68
	(b"10111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111011000010100011110101110", b"10111111100010111000010100011111"), -- -0.21 + -0.88 = -1.09
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111110001110000101000111101100", b"00111111010000000000000000000000"), -- 0.57 + 0.18 = 0.75
	(b"00111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"00111111100000101000111101011100"), -- 0.03 + 0.99 = 1.02
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111011110000101000111101100"), -- -0.17 + -0.8 = -0.97
	(b"10111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111001100110011001100110011"), -- -0.12 + -0.58 = -0.7
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011100110011001100110011", b"00111111011111010111000010100100"), -- 0.04 + 0.95 = 0.99
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"10111111111010100011110101110000"), -- -0.87 + -0.96 = -1.83
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"10111111101100011110101110000110"), -- -0.54 + -0.85 = -1.39
	(b"10111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000111000010100011110110"), -- -0.11 + -0.5 = -0.61
	(b"00111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111111010101000111101011100001"), -- 0.75 + 0.08 = 0.83
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111110001010001111010111000"), -- -0.64 + -0.9 = -1.54
	(b"00111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111111100011110101110000101001"), -- 0.33 + 0.79 = 1.12
	(b"00111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111001100110011001100110011"), -- 0.46 + 0.24 = 0.7
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111001110000101000111101100", b"10111111110001111010111000010100"), -- -0.84 + -0.72 = -1.56
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"00111111110111010111000010100100"), -- 0.86 + 0.87 = 1.73
	(b"10111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111111010100011110101110000101"), -- -0.44 + -0.38 = -0.82
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"00111111011100110011001100110011"), -- 0.7 + 0.25 = 0.95
	(b"10111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001110000101000111101100", b"10111111110101011100001010010000"), -- -0.95 + -0.72 = -1.67
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111100111000010100011110110"), -- -0.79 + -0.43 = -1.22
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001001100110011001100110", b"10111111110011100001010001111010"), -- -0.96 + -0.65 = -1.61
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111101101000111101011100010"), -- -0.61 + -0.8 = -1.41
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111100000111101011100001010"), -- -0.09 + -0.94 = -1.03
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111100100110011001100110011"), -- 0.63 + 0.52 = 1.15
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111101111010111000010100100"), -- -0.79 + -0.69 = -1.48
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111100100001010001111010111"), -- 0.37 + 0.76 = 1.13
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"10111111100100001010001111010111"), -- -0.24 + -0.89 = -1.13
	(b"10111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111000011001100110011001101", b"10111111101101110000101000111110"), -- -0.88 + -0.55 = -1.43
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111111100000101000111101011100"), -- 0.97 + 0.05 = 1.02
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"00111111011000111101011100001010"), -- 0.56 + 0.33 = 0.89
	(b"00111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"00111111101010100011110101110000"), -- 0.94 + 0.39 = 1.33
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111010010100011110101110001"), -- -0.79 + -0 = -0.79
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111010101110000101000111110"), -- -0.23 + -0.61 = -0.84
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"10111111000011110101110000101001"), -- -0.3 + -0.26 = -0.56
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110000001010001111010111000", b"10111111000101000111101011100001"), -- -0.45 + -0.13 = -0.58
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111110110101110000101001000"), -- 0.95 + 0.76 = 1.71
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111001111010111000010100100"), -- -0.17 + -0.57 = -0.74
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111011110000101000111101100", b"10111111100110011001100110011010"), -- -0.23 + -0.97 = -1.2
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"00111111101000101000111101011100"), -- 0.43 + 0.84 = 1.27
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111011000010100011110101110", b"10111111100011110101110000101001"), -- -0.24 + -0.88 = -1.12
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111100000101000111101011100"), -- -0.4 + -0.62 = -1.02
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"10111111100100110011001100110011"), -- -0.4 + -0.75 = -1.15
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111110110001111010111000010100"), -- 0.01 + 0.38 = 0.39
	(b"10111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110000110011001100110011010", b"10111111000000000000000000000000"), -- -0.35 + -0.15 = -0.5
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111011001100110011001100111"), -- 0.36 + 0.54 = 0.9
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111010001010001111010111000", b"00111111110100001010001111010111"), -- 0.86 + 0.77 = 1.63
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111101001010001111010111000"), -- -0.72 + -0.57 = -1.29
	(b"10111110100111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111011011100001010001111011"), -- -0.31 + -0.62 = -0.93
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111010111000010100011110101"), -- 0.21 + 0.65 = 0.86
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110101000111101011100001010", b"00111110101011100001010001111011"), -- 0.02 + 0.32 = 0.34
	(b"00111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111100110011001100110011010"), -- 0.53 + 0.67 = 1.2
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111101000111101011100001010"), -- 0.4 + 0.88 = 1.28
	(b"00111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111100100110011001100110011"), -- 0.51 + 0.64 = 1.15
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111110100110011001100110011"), -- 0.89 + 0.76 = 1.65
	(b"00111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111111100101110000101000111110"), -- 0.75 + 0.43 = 1.18
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111110100110011001100110011"), -- 0.95 + 0.7 = 1.65
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111110011001100110011001100"), -- -0.9 + -0.7 = -1.6
	(b"10111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"10111111100000010100011110101110"), -- -0.85 + -0.16 = -1.01
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010100011110101110000101", b"00111111111000101000111101011100"), -- 0.95 + 0.82 = 1.77
	(b"00111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111011101011100001010001111", b"00111111101011110101110000101001"), -- 0.41 + 0.96 = 1.37
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111101000101000111101011100"), -- 0.62 + 0.65 = 1.27
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010001010001111010111000", b"00111111110111000010100011110110"), -- 0.95 + 0.77 = 1.72
	(b"10111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"10111111101111000010100011110110"), -- -0.73 + -0.74 = -1.47
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111111100110101110000101001000"), -- -0.76 + -0.45 = -1.21
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111101010100011110101110000"), -- -0.53 + -0.8 = -1.33
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111101101110000101000111101100", b"00111111001000010100011110101110"), -- 0.54 + 0.09 = 0.63
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111110111101011100001010010"), -- -0.9 + -0.84 = -1.74
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111001101011100001010001111", b"10111111010101110000101000111101"), -- -0.13 + -0.71 = -0.84
	(b"10111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111100110011001100110011010"), -- -0.59 + -0.61 = -1.2
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111101000010100011110101110"), -- 0.62 + 0.64 = 1.26
	(b"00111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111111100110101110000101001000"), -- 0.83 + 0.38 = 1.21
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111001010001111010111000011", b"10111111010010100011110101110001"), -- -0.13 + -0.66 = -0.79
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111000000000000000000000000"), -- -0.09 + -0.41 = -0.5
	(b"10111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111100101011100001010001111"), -- -0.59 + -0.58 = -1.17
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111100011001100110011001101"), -- -0.77 + -0.33 = -1.1
	(b"00111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"00111111000001010001111010111000"), -- 0.46 + 0.06 = 0.52
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110111110101110000101001000", b"10111111100101000111101011100010"), -- -0.67 + -0.49 = -1.16
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011110000101000111101100", b"10111111100101011100001010010000"), -- -0.2 + -0.97 = -1.17
	(b"10111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111111011110101110000101001"), -- -0.97 + -0.9 = -1.87
	(b"00111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111111010000101000111101011100"), -- 0.71 + 0.05 = 0.76
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111111100100001010001111010111"), -- 0.97 + 0.16 = 1.13
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111001010001111010111000011", b"10111111011100001010001111011000"), -- -0.28 + -0.66 = -0.94
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"10111111100110011001100110011010"), -- -0.76 + -0.44 = -1.2
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"00111110110100011110101110000101"), -- 0.34 + 0.07 = 0.41
	(b"00111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110110100011110101110000101", b"00111111000001111010111000010100"), -- 0.12 + 0.41 = 0.53
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110100010100011110101110001", b"00111110111000010100011110101110"), -- 0.17 + 0.27 = 0.44
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"00111111100000000000000000000000"), -- 0.97 + 0.03 = 1
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111100100110011001100110011"), -- -0.45 + -0.7 = -1.15
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001011100001010001111011", b"00111111100101110000101000111110"), -- 0.5 + 0.68 = 1.18
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111101111101011100001010001111", b"00111110101110000101000111101011"), -- 0.24 + 0.12 = 0.36
	(b"00111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111010101000111101011100001"), -- 0.19 + 0.64 = 0.83
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111101100110011001100110011"), -- 0.59 + 0.81 = 1.4
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111101010100011110101110000"), -- -0.71 + -0.62 = -1.33
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111011110101110000101001000", b"10111111100011100001010001111011"), -- -0.13 + -0.98 = -1.11
	(b"00111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111100000000000000000000000"), -- 0.51 + 0.49 = 1
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111111011001100110011001100"), -- 0.95 + 0.9 = 1.85
	(b"10111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"10111111101010100011110101110000"), -- -0.59 + -0.74 = -1.33
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110111010111000010100011111", b"10111111100101110000101000111110"), -- -0.72 + -0.46 = -1.18
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111001010111000010100011111"), -- -0.05 + -0.62 = -0.67
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111101001100110011001100110"), -- 0.6 + 0.7 = 1.3
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111100100001010001111010111"), -- 0.73 + 0.4 = 1.13
	(b"00111111011011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111110110000101000111101100"), -- 0.93 + 0.76 = 1.69
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111100000111101011100001010"), -- 0.57 + 0.46 = 1.03
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010011110101110000101001", b"10111111100001010001111010111000"), -- -0.23 + -0.81 = -1.04
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110101111010111000010100100", b"10111111100101011100001010010000"), -- -0.8 + -0.37 = -1.17
	(b"10111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111100100001010001111010111"), -- -0.56 + -0.57 = -1.13
	(b"00111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110100010100011110101110001", b"00111111100011001100110011001101"), -- 0.83 + 0.27 = 1.1
	(b"00111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111100001010001111010111000"), -- 0.58 + 0.46 = 1.04
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"00111111000110011001100110011010"), -- 0.29 + 0.31 = 0.6
	(b"10111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110110101110000101000111101", b"10111111001000010100011110101110"), -- -0.21 + -0.42 = -0.63
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000001111010111000010100", b"00111111000101000111101011100001"), -- 0.05 + 0.53 = 0.58
	(b"00111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111111010001010001111010111000"), -- 0.28 + 0.49 = 0.77
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011101011100001010001111", b"00111111111000010100011110101110"), -- 0.8 + 0.96 = 1.76
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111111011100001010001111010111"), -- 0.81 + 0.13 = 0.94
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111100010111000010100011111"), -- -0.48 + -0.61 = -1.09
	(b"00111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111110111100001010001111011000"), -- 0.33 + 0.14 = 0.47
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110101100110011001100110011", b"10111111010001010001111010111000"), -- -0.42 + -0.35 = -0.77
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"10111111111100001010001111010111"), -- -0.92 + -0.96 = -1.88
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001101011100001010001111", b"00111111101001111010111000010100"), -- 0.6 + 0.71 = 1.31
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111100011110101110000101001"), -- 0.78 + 0.34 = 1.12
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111110011110101110000101001"), -- 0.73 + 0.89 = 1.62
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"00111111100001111010111000010100"), -- 0.59 + 0.47 = 1.06
	(b"00111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011010111000010100011111", b"00111111111100001010001111010111"), -- 0.96 + 0.92 = 1.88
	(b"00111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111101111101011100001010001111", b"00111111100001010001111010111000"), -- 0.92 + 0.12 = 1.04
	(b"00111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111010011110101110000101001", b"00111111101111000010100011110110"), -- 0.66 + 0.81 = 1.47
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111011110000101000111101100", b"10111111101011100001010001111011"), -- -0.39 + -0.97 = -1.36
	(b"10111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111011100110011001100110011"), -- -0.44 + -0.51 = -0.95
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"00111111110011110101110000101001"), -- 0.97 + 0.65 = 1.62
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"00111111010101110000101000111110"), -- 0.56 + 0.28 = 0.84
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111100110101110000101001000"), -- 0.32 + 0.89 = 1.21
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111111101000111101011100001010"), -- -0.83 + -0.45 = -1.28
	(b"00111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111100101000111101011100001"), -- 0.64 + 0.52 = 1.16
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111100011110101110000101001"), -- 0.78 + 0.34 = 1.12
	(b"00111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111110111001100110011001100110"), -- 0.07 + 0.38 = 0.45
	(b"10111110111100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"10111111101001010001111010111000"), -- -0.47 + -0.82 = -1.29
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111101011101011100001010001111", b"10111111001010111000010100011111"), -- -0.61 + -0.06 = -0.67
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111111011001100110011001101"), -- -0.86 + -0.99 = -1.85
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111110111010111000010100100"), -- -0.79 + -0.94 = -1.73
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111011000111101011100001010"), -- 0.22 + 0.67 = 0.89
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"00111111001110000101000111101011"), -- 0.69 + 0.03 = 0.72
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110100011110101110000101001", b"10111110110100011110101110000101"), -- -0.13 + -0.28 = -0.41
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111001010111000010100011111"), -- -0.36 + -0.31 = -0.67
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111010000101000111101011100"), -- 0.24 + 0.52 = 0.76
	(b"00111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111010110011001100110011010", b"00111111011101011100001010010000"), -- 0.11 + 0.85 = 0.96
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"10111111010010100011110101110000"), -- -0.78 + -0.01 = -0.79
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"10111111101010001111010111000010"), -- -0.43 + -0.89 = -1.32
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111010000101000111101011100", b"10111111101000000000000000000000"), -- -0.49 + -0.76 = -1.25
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111100100001010001111010111"), -- -0.52 + -0.61 = -1.13
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111001011100001010001111011", b"10111111100010100011110101110001"), -- -0.4 + -0.68 = -1.08
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111100111010111000010100100"), -- -0.54 + -0.69 = -1.23
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000101000111101011100", b"00111111100001111010111000010100"), -- 0.55 + 0.51 = 1.06
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111001010111000010100011111", b"10111111101110000101000111101100"), -- -0.77 + -0.67 = -1.44
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111100001010001111010111000"), -- -0.2 + -0.84 = -1.04
	(b"00111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"00111111100000000000000000000000"), -- 0.45 + 0.55 = 1
	(b"10111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111101011001100110011001100"), -- -0.51 + -0.84 = -1.35
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111101011100001010001111011"), -- 0.86 + 0.5 = 1.36
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"10111111101011001100110011001101"), -- -0.36 + -0.99 = -1.35
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"00111111010010100011110101110001"), -- 0.62 + 0.17 = 0.79
	(b"00111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011011100001010001111011", b"00111111100010100011110101110001"), -- 0.15 + 0.93 = 1.08
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"00111110111010111000010100011110"), -- 0.01 + 0.45 = 0.46
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111111010100011110101110000101"), -- 0.74 + 0.08 = 0.82
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101111000010100011110101110", b"00111110101110000101000111101100"), -- 0.25 + 0.11 = 0.36
	(b"00111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111101001010001111010111000"), -- 0.46 + 0.83 = 1.29
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111001000111101011100001010", b"00111111101001111010111000010100"), -- 0.67 + 0.64 = 1.31
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"10111111010111000010100011110110"), -- -0.01 + -0.85 = -0.86
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110001111010111000010100", b"10111111010101110000101000111101"), -- -0.45 + -0.39 = -0.84
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111010101110000101000111110"), -- 0.3 + 0.54 = 0.84
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111110001110000101000111101100"), -- 0.04 + 0.14 = 0.18
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111011100001010001111010111"), -- -0.24 + -0.7 = -0.94
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111110101000111101011100001"), -- -0.71 + -0.95 = -1.66
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111000011001100110011001101"), -- -0.24 + -0.31 = -0.55
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111001101011100001010001111", b"00111111100010001111010111000010"), -- 0.36 + 0.71 = 1.07
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110010101110000101000111101", b"00111111000011001100110011001101"), -- 0.34 + 0.21 = 0.55
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111110010001111010111000010"), -- 0.69 + 0.88 = 1.57
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011110101110000101001000", b"00111111110000111101011100001010"), -- 0.55 + 0.98 = 1.53
	(b"00111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111001000010100011110101110", b"00111111101110011001100110011010"), -- 0.82 + 0.63 = 1.45
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111011101011100001010001111"), -- -0.01 + -0.95 = -0.96
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111101110101110000101001000"), -- 0.63 + 0.83 = 1.46
	(b"00111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111100001000111101011100001010", b"00111111010101000111101011100001"), -- 0.82 + 0.01 = 0.83
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111100001111010111000010100"), -- -0.45 + -0.61 = -1.06
	(b"00111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111001110101110000101001000"), -- 0.39 + 0.34 = 0.73
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111110101111010111000010100100", b"10111111010111000010100011110110"), -- -0.49 + -0.37 = -0.86
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011010001111010111000011", b"10111111100000010100011110101110"), -- -0.1 + -0.91 = -1.01
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111000001111010111000010100"), -- -0 + -0.53 = -0.53
	(b"00111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111100111010111000010100100"), -- 0.71 + 0.52 = 1.23
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111001010001111010111000010"), -- -0.13 + -0.53 = -0.66
	(b"00111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111101100001010001111010111"), -- 0.62 + 0.76 = 1.38
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110101011100001010001111011", b"10111111010111101011100001010010"), -- -0.53 + -0.34 = -0.87
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111001011100001010001111011", b"00111111100110011001100110011010"), -- 0.52 + 0.68 = 1.2
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111101101011100001010010000"), -- -0.72 + -0.7 = -1.42
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111101110011001100110011010"), -- -0.92 + -0.53 = -1.45
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111110110111000010100011110110"), -- 0.35 + 0.08 = 0.43
	(b"10111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"10111111100100110011001100110011"), -- -0.41 + -0.74 = -1.15
	(b"00111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"00111111111001010001111010111000"), -- 0.85 + 0.94 = 1.79
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001011100001010001111011", b"00111111010001111010111000010101"), -- 0.1 + 0.68 = 0.78
	(b"00111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"00111111010101000111101011100001"), -- 0.77 + 0.06 = 0.83
	(b"10111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111011010001111010111000010"), -- -0.32 + -0.59 = -0.91
	(b"10111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111010001010001111010111000", b"10111111101000111101011100001010"), -- -0.51 + -0.77 = -1.28
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111011010001111010111000011", b"00111111110011001100110011001101"), -- 0.69 + 0.91 = 1.6
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111110000111101011100001010"), -- -0.69 + -0.84 = -1.53
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"10111110010101110000101000111101"), -- -0.13 + -0.08 = -0.21
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111101001100110011001100110"), -- -0.43 + -0.87 = -1.3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"00111111101001010001111010111000"), -- 0.9 + 0.39 = 1.29
	(b"10111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111101101110000101000111101100", b"10111110110100011110101110000101"), -- -0.32 + -0.09 = -0.41
	(b"00111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111110011001100110011001100"), -- 0.71 + 0.89 = 1.6
	(b"00111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111001111010111000010100100", b"00111111011000010100011110101110"), -- 0.14 + 0.74 = 0.88
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000001010001111010111000", b"10111111000101000111101011100001"), -- -0.06 + -0.52 = -0.58
	(b"10111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111110110100011110101110000101"), -- -0.41 + -0 = -0.41
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"00111111100000000000000000000000"), -- 0.78 + 0.22 = 1
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111111010001010001111010111001"), -- 0.72 + 0.05 = 0.77
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011110101110000101001000", b"10111111100101110000101000111110"), -- -0.2 + -0.98 = -1.18
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111001110000101000111101100", b"10111111101100011110101110000110"), -- -0.67 + -0.72 = -1.39
	(b"10111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"10111111001111010111000010100100"), -- -0.62 + -0.12 = -0.74
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111011011100001010001111011"), -- 0.73 + 0.2 = 0.93
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111100010111000010100011111"), -- 0.63 + 0.46 = 1.09
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111111010110011001100110011010"), -- 0.69 + 0.16 = 0.85
	(b"10111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111101110101110000101001000"), -- -0.67 + -0.79 = -1.46
	(b"00111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111001111010111000010100100", b"00111111110000000000000000000000"), -- 0.76 + 0.74 = 1.5
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"10111111001000010100011110101110"), -- -0.45 + -0.18 = -0.63
	(b"10111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111010111000010100011110110", b"10111111101101011100001010010000"), -- -0.56 + -0.86 = -1.42
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111001000010100011110101110"), -- 0.29 + 0.34 = 0.63
	(b"10111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"10111111100100001010001111010111"), -- -0.91 + -0.22 = -1.13
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111100000111101011100001010"), -- 0.3 + 0.73 = 1.03
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111011100110011001100110011"), -- 0.43 + 0.52 = 0.95
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"10111111101001100110011001100110"), -- -0.86 + -0.44 = -1.3
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"10111111100011100001010001111011"), -- -0.15 + -0.96 = -1.11
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111111010111000010100011110"), -- -0.89 + -0.95 = -1.84
	(b"00111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"00111111101000101000111101011100"), -- 0.98 + 0.29 = 1.27
	(b"10111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111110100110011001100110100"), -- -0.85 + -0.8 = -1.65
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"10111111001110000101000111101011"), -- -0.69 + -0.03 = -0.72
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111001111010111000010100100"), -- -0.24 + -0.5 = -0.74
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111010011110101110000101001", b"10111111101101011100001010010000"), -- -0.61 + -0.81 = -1.42
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111111011001100110011001100110"), -- -0.52 + -0.38 = -0.9
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110101000111101011100001010", b"10111111100000101000111101011100"), -- -0.7 + -0.32 = -1.02
	(b"00111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111101101110000101000111101100", b"00111110101010001111010111000010"), -- 0.24 + 0.09 = 0.33
	(b"00111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"00111111000001010001111010111000"), -- 0.13 + 0.39 = 0.52
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"10111111101010100011110101110000"), -- -0.37 + -0.96 = -1.33
	(b"10111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111111100001111010111000010100"), -- -0.68 + -0.38 = -1.06
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110101000111101011100001010", b"10111111100011100001010001111011"), -- -0.79 + -0.32 = -1.11
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111101100110011001100110011"), -- -0.89 + -0.51 = -1.4
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111011100001010001111010111"), -- -0.3 + -0.64 = -0.94
	(b"00111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111111101011110101110000101001"), -- 0.99 + 0.38 = 1.37
	(b"00111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"00111111100011110101110000101001"), -- 0.28 + 0.84 = 1.12
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"10111111100001111010111000010100"), -- -0.23 + -0.83 = -1.06
	(b"10111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111111000110011001100110011010"), -- -0.22 + -0.38 = -0.6
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111010100011110101110000101", b"00111111100110011001100110011010"), -- 0.38 + 0.82 = 1.2
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"00111111110001111010111000010100"), -- 0.59 + 0.97 = 1.56
	(b"00111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"00111110110000101000111101011100"), -- 0.07 + 0.31 = 0.38
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000111000010100011110110", b"00111111100011100001010001111011"), -- 0.5 + 0.61 = 1.11
	(b"10111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111001010001111010111000010"), -- -0.13 + -0.53 = -0.66
	(b"00111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"00111111100011110101110000101001"), -- 0.15 + 0.97 = 1.12
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010110011001100110011010", b"00111111111001100110011001100110"), -- 0.95 + 0.85 = 1.8
	(b"00111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"00111111101101110000101000111110"), -- 0.88 + 0.55 = 1.43
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"00111111100010100011110101110001"), -- 0.79 + 0.29 = 1.08
	(b"10111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"10111111111000010100011110101110"), -- -0.94 + -0.82 = -1.76
	(b"00111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"00111101111000010100011110101110"), -- 0.06 + 0.05 = 0.11
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010010100011110101110001", b"10111111011111010111000010100100"), -- -0.2 + -0.79 = -0.99
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"10111111000001111010111000010100"), -- -0.52 + -0.01 = -0.53
	(b"00111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"00111111110111010111000010100100"), -- 0.76 + 0.97 = 1.73
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111011100110011001100110011", b"00111111100101011100001010001111"), -- 0.22 + 0.95 = 1.17
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111100001111010111000010100"), -- 0.23 + 0.83 = 1.06
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"10111111101101110000101000111110"), -- -0.69 + -0.74 = -1.43
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"00111111010111000010100011110110"), -- 0.55 + 0.31 = 0.86
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111011000111101011100001010"), -- -0.36 + -0.53 = -0.89
	(b"00111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111100111000010100011110110"), -- 0.98 + 0.24 = 1.22
	(b"00111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"00111110101110000101000111101100"), -- 0.19 + 0.17 = 0.36
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111110110100011110101110000101"), -- -0.39 + -0.02 = -0.41
	(b"00111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111100101000111101011100010"), -- 0.49 + 0.67 = 1.16
	(b"00111110111100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111001101011100001010001111"), -- 0.47 + 0.24 = 0.71
	(b"10111110100111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111010101110000101000111101"), -- -0.31 + -0.53 = -0.84
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111010101110000101000111110"), -- 0.3 + 0.54 = 0.84
	(b"00111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111011010001111010111000010"), -- 0.57 + 0.34 = 0.91
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"00111111001110000101000111101100"), -- 0.35 + 0.37 = 0.72
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"00111111000011110101110000101001"), -- 0.04 + 0.52 = 0.56
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110110111000010100011110110", b"00111110111001100110011001100111"), -- 0.02 + 0.43 = 0.45
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110110101110000101000111101", b"00111110110111000010100011110101"), -- 0.01 + 0.42 = 0.43
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111100110101110000101001000"), -- -0.78 + -0.43 = -1.21
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110001111010111000010100", b"10111111001100001010001111010111"), -- -0.3 + -0.39 = -0.69
	(b"10111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011000010100011110101110", b"10111111011001100110011001100110"), -- -0.02 + -0.88 = -0.9
	(b"00111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111011110101110000101001000", b"00111111100101011100001010010000"), -- 0.19 + 0.98 = 1.17
	(b"00111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111001111010111000010100100", b"00111111100100110011001100110011"), -- 0.41 + 0.74 = 1.15
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"00111111000110011001100110011010"), -- 0.56 + 0.04 = 0.6
	(b"10111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111101000010100011110101110"), -- -0.75 + -0.51 = -1.26
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"10111111011110101110000101001000"), -- -0.8 + -0.18 = -0.98
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001011100001010001111011", b"10111111101100011110101110000101"), -- -0.71 + -0.68 = -1.39
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111101001111010111000010101"), -- 0.97 + 0.34 = 1.31
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111101111000010100011110101110", b"00111111010101000111101011100010"), -- 0.72 + 0.11 = 0.83
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"00111110101010001111010111000011"), -- 0.05 + 0.28 = 0.33
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"10111111110100110011001100110011"), -- -0.82 + -0.83 = -1.65
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110111000010100011110101110", b"00111110111010111000010100011111"), -- 0.02 + 0.44 = 0.46
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111010011001100110011001101"), -- 0.04 + 0.76 = 0.8
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110011000010100011110101110", b"10111111100011100001010001111011"), -- -0.89 + -0.22 = -1.11
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"10111110010101110000101000111110"), -- -0.04 + -0.17 = -0.21
	(b"10111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111000101000111101011100010"), -- -0.15 + -0.43 = -0.58
	(b"00111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111000010100011110101110001"), -- 0.14 + 0.4 = 0.54
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111100010001111010111000010"), -- 0.17 + 0.9 = 1.07
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"10111111101010100011110101110000"), -- -0.71 + -0.62 = -1.33
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111111000000000000000000000000"), -- 0.36 + 0.14 = 0.5
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110011010111000010100011111", b"00111111000101000111101011100001"), -- 0.35 + 0.23 = 0.58
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110101000111101011100001010", b"10111111001111010111000010100100"), -- -0.42 + -0.32 = -0.74
	(b"10111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"10111111100000000000000000000000"), -- -0.99 + -0.01 = -1
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111111100101011100001010010000"), -- 0.55 + 0.62 = 1.17
	(b"00111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110100010100011110101110001", b"00111111100110101110000101001000"), -- 0.94 + 0.27 = 1.21
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011010111000010100011111", b"10111111100111000010100011110110"), -- -0.3 + -0.92 = -1.22
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111101000000000000000000000"), -- -0.84 + -0.41 = -1.25
	(b"10111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111110100001010001111010111000"), -- -0.07 + -0.19 = -0.26
	(b"10111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111001010001111010111000011", b"10111111101010111000010100011111"), -- -0.68 + -0.66 = -1.34
	(b"00111110000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111110000110011001100110011010"), -- 0.15 + 0 = 0.15
	(b"10111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111010000000000000000000000"), -- -0.22 + -0.53 = -0.75
	(b"10111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111101011110101110000101001"), -- -0.74 + -0.63 = -1.37
	(b"00111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"00111111001000111101011100001010"), -- 0.33 + 0.31 = 0.64
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111110101111010111000010100100"), -- 0.21 + 0.16 = 0.37
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010101110000101000111101", b"00111110110100011110101110000101"), -- 0.2 + 0.21 = 0.41
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100010100011110101110001", b"10111111001010111000010100011111"), -- -0.4 + -0.27 = -0.67
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111010001111010111000010100", b"00111111110000101000111101011100"), -- 0.74 + 0.78 = 1.52
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"10111111110011001100110011001100"), -- -0.77 + -0.83 = -1.6
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"10111110111010111000010100011110"), -- -0.45 + -0.01 = -0.46
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111001110101110000101001000", b"00111111100010111000010100011111"), -- 0.36 + 0.73 = 1.09
	(b"10111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111011000111101011100001010"), -- -0.19 + -0.7 = -0.89
	(b"00111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"00111111011100001010001111010111"), -- 0.07 + 0.87 = 0.94
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111010110011001100110011010"), -- -0.24 + -0.61 = -0.85
	(b"00111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"00111111100010111000010100011111"), -- 0.87 + 0.22 = 1.09
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111101110000101000111101100"), -- 0.86 + 0.58 = 1.44
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110100010100011110101110001", b"10111111001000010100011110101110"), -- -0.36 + -0.27 = -0.63
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110100101000111101011100001", b"10111111000001111010111000010100"), -- -0.24 + -0.29 = -0.53
	(b"00111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110101011100001010001111011", b"00111111010001111010111000010100"), -- 0.44 + 0.34 = 0.78
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"00111110111110101110000101001000"), -- 0.3 + 0.19 = 0.49
	(b"10111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110110001111010111000010100"), -- -0.19 + -0.2 = -0.39
	(b"10111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110101011100001010001111011", b"10111111011001100110011001100110"), -- -0.56 + -0.34 = -0.9
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111010110011001100110011010"), -- -0.52 + -0.33 = -0.85
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111111001010111000010100011110"), -- 0.29 + 0.38 = 0.67
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"10111111001110101110000101001000"), -- -0.4 + -0.33 = -0.73
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"10111110100011110101110000101001"), -- -0.2 + -0.08 = -0.28
	(b"10111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111010011001100110011001101"), -- -0.11 + -0.69 = -0.8
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"00111110100001010001111010111000"), -- 0.1 + 0.16 = 0.26
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111110000010100011110101110"), -- -0.81 + -0.7 = -1.51
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000001010001111010111000", b"10111111011110000101000111101011"), -- -0.45 + -0.52 = -0.97
	(b"10111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"10111111011000010100011110101110"), -- -0.35 + -0.53 = -0.88
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"10111111100100011110101110000101"), -- -0.36 + -0.78 = -1.14
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111100101000111101011100001010", b"10111111000111101011100001010010"), -- -0.6 + -0.02 = -0.62
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111101111101011100001010010"), -- 0.95 + 0.54 = 1.49
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"10111110101010001111010111000010"), -- -0.16 + -0.17 = -0.33
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111110000000000000000000000"), -- -0.87 + -0.63 = -1.5
	(b"10111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111111001010001111010111000"), -- -0.85 + -0.94 = -1.79
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111111010111000010100011110"), -- -0.9 + -0.94 = -1.84
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"10111111100010100011110101110000"), -- -0.3 + -0.78 = -1.08
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011010001111010111000011", b"00111111101101000111101011100010"), -- 0.5 + 0.91 = 1.41
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111001011100001010001111011", b"00111111101011001100110011001101"), -- 0.67 + 0.68 = 1.35
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111100100110011001100110011"), -- -0.25 + -0.9 = -1.15
	(b"10111111000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"10111111101001111010111000010100"), -- -0.62 + -0.69 = -1.31
	(b"00111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111110111000010100011110101110", b"00111111010101000111101011100001"), -- 0.39 + 0.44 = 0.83
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"00111111100000101000111101011100"), -- 0.8 + 0.22 = 1.02
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110110101110000101000111101", b"10111111100001111010111000010100"), -- -0.64 + -0.42 = -1.06
	(b"10111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"10111111100010001111010111000011"), -- -0.99 + -0.08 = -1.07
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110010101110000101000111101", b"10111110111000010100011110101110"), -- -0.23 + -0.21 = -0.44
	(b"00111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111000100011110101110000101"), -- 0.33 + 0.24 = 0.57
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111100011001100110011001101"), -- -0.16 + -0.94 = -1.1
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111001110000101000111101100", b"00111111110000010100011110101110"), -- 0.79 + 0.72 = 1.51
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"10111111010001111010111000010100"), -- -0.14 + -0.64 = -0.78
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110010101110000101000111101", b"00111110011010111000010100011110"), -- 0.02 + 0.21 = 0.23
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111100100011110101110000101"), -- -0.84 + -0.3 = -1.14
	(b"00111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"00111111001000010100011110101110"), -- 0.26 + 0.37 = 0.63
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"00111111011010111000010100011110"), -- 0.59 + 0.33 = 0.92
	(b"00111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"00111111101011110101110000101000"), -- 0.53 + 0.84 = 1.37
	(b"10111110100111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"10111111101000000000000000000000"), -- -0.31 + -0.94 = -1.25
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"00111111100111000010100011110110"), -- 0.35 + 0.87 = 1.22
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111010111101011100001010010", b"10111111101101000111101011100010"), -- -0.54 + -0.87 = -1.41
	(b"00111111011011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110000011110101110000101001", b"00111111100010001111010111000011"), -- 0.93 + 0.14 = 1.07
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111001010001111010111000011", b"00111111010111101011100001010010"), -- 0.21 + 0.66 = 0.87
	(b"00111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"00111111100110000101000111101100"), -- 0.65 + 0.54 = 1.19
	(b"10111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110110001111010111000010100", b"10111111000101000111101011100001"), -- -0.19 + -0.39 = -0.58
	(b"10111101100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111011010001111010111000010"), -- -0.07 + -0.84 = -0.91
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111101100110011001100110011"), -- -0.83 + -0.57 = -1.4
	(b"00111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111101010111000010100011110"), -- 0.76 + 0.58 = 1.34
	(b"10111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111010111000010100011110110"), -- -0.66 + -0.2 = -0.86
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"00111111100111101011100001010010"), -- 0.79 + 0.45 = 1.24
	(b"10111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011010111000010100011111", b"10111111111000101000111101011100"), -- -0.85 + -0.92 = -1.77
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"10111111100101011100001010010000"), -- -0.43 + -0.74 = -1.17
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010110011001100110011010", b"00111111110100110011001100110100"), -- 0.8 + 0.85 = 1.65
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111100001111010111000010100"), -- 0.23 + 0.83 = 1.06
	(b"00111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"00111110010000101000111101011100"), -- 0.16 + 0.03 = 0.19
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111001110101110000101001000", b"10111111101011110101110000101001"), -- -0.64 + -0.73 = -1.37
	(b"00111101111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"00111110010000101000111101011100"), -- 0.12 + 0.07 = 0.19
	(b"00111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111011110101110000101001000"), -- 0.09 + 0.89 = 0.98
	(b"10111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110011101011100001010001111", b"10111111010000000000000000000000"), -- -0.51 + -0.24 = -0.75
	(b"10111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111111011100001010001111010111"), -- -0.75 + -0.19 = -0.94
	(b"00111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111100101000111101011100001"), -- 0.96 + 0.2 = 1.16
	(b"10111111001101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111010011110101110000101001"), -- -0.71 + -0.1 = -0.81
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111100001100110011001100110"), -- -0.64 + -0.41 = -1.05
	(b"10111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"10111111011100001010001111010111"), -- -0.91 + -0.03 = -0.94
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"00111111100011001100110011001100"), -- 0.52 + 0.58 = 1.1
	(b"00111111001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111000100011110101110000101", b"00111111100111101011100001010010"), -- 0.67 + 0.57 = 1.24
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111110100101000111101011100001"), -- 0.21 + 0.08 = 0.29
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"00111111100100011110101110000101"), -- 0.9 + 0.24 = 1.14
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110100111101011100001010010", b"10111111100000010100011110101110"), -- -0.7 + -0.31 = -1.01
	(b"10111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"10111111001010111000010100011111"), -- -0.55 + -0.12 = -0.67
	(b"10111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110010101110000101000111101", b"10111111000101110000101000111101"), -- -0.38 + -0.21 = -0.59
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110101110000101000111101100", b"00111111100101011100001010010000"), -- 0.81 + 0.36 = 1.17
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111101101110000101000111110"), -- 0.6 + 0.83 = 1.43
	(b"10111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"10111111001001100110011001100110"), -- -0.46 + -0.19 = -0.65
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111001000010100011110101110", b"10111111100001100110011001100110"), -- -0.42 + -0.63 = -1.05
	(b"10111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111000111000010100011110110", b"10111111100101110000101000111110"), -- -0.57 + -0.61 = -1.18
	(b"00111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"00111111100000010100011110101110"), -- 0.04 + 0.97 = 1.01
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"00111111000010100011110101110001"), -- 0.5 + 0.04 = 0.54
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"00111111011000111101011100001010"), -- 0.5 + 0.39 = 0.89
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"00111111100000111101011100001010"), -- 0.95 + 0.08 = 1.03
	(b"00111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011011100001010001111011", b"00111111110101110000101000111110"), -- 0.75 + 0.93 = 1.68
	(b"10111110010000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"10111110101100110011001100110011"), -- -0.19 + -0.16 = -0.35
	(b"00111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00111110001011100001010001111011"), -- 0.17 + 0 = 0.17
	(b"00111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111000011110101110000101001", b"00111111101101011100001010010000"), -- 0.86 + 0.56 = 1.42
	(b"00111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111001101011100001010001111", b"00111111110011110101110000101001"), -- 0.91 + 0.71 = 1.62
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"10111111101100011110101110000101"), -- -0.5 + -0.89 = -1.39
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110010000101000111101011100", b"00111111100010111000010100011110"), -- 0.9 + 0.19 = 1.09
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110111101011100001010001111", b"10111111001011100001010001111011"), -- -0.2 + -0.48 = -0.68
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111100110011001100110011010"), -- 0.5 + 0.7 = 1.2
	(b"10111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111011011100001010001111011", b"10111111110011100001010001111011"), -- -0.68 + -0.93 = -1.61
	(b"10111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110100010100011110101110001", b"10111111000101110000101000111110"), -- -0.32 + -0.27 = -0.59
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110101100110011001100110011", b"00111110101100110011001100110011"), -- 0 + 0.35 = 0.35
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111100000111101011100001010"), -- 0.63 + 0.4 = 1.03
	(b"10111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"10111111000110011001100110011001"), -- -0.02 + -0.58 = -0.6
	(b"10111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111110001100110011001100110"), -- -0.75 + -0.8 = -1.55
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"10111111100100110011001100110011"), -- -0.37 + -0.78 = -1.15
	(b"00111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111000000101000111101011100", b"00111111000110011001100110011010"), -- 0.09 + 0.51 = 0.6
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"10111101101110000101000111101100"), -- -0.05 + -0.04 = -0.09
	(b"00111111011010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111010000101000111101011100", b"00111111110101011100001010010000"), -- 0.91 + 0.76 = 1.67
	(b"00111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110101111010111000010100100", b"00111110110011001100110011001101"), -- 0.03 + 0.37 = 0.4
	(b"00111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010000000000000000000000", b"00111111010001010001111010111000"), -- 0.02 + 0.75 = 0.77
	(b"00111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011010111000010100011111", b"00111111100000000000000000000000"), -- 0.08 + 0.92 = 1
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010111101011100001010010", b"00111111011000010100011110101110"), -- 0.01 + 0.87 = 0.88
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"00111110110111000010100011110110"), -- 0.05 + 0.38 = 0.43
	(b"00111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"00111111101000101000111101011100"), -- 0.48 + 0.79 = 1.27
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"00111111010000000000000000000000"), -- 0.72 + 0.03 = 0.75
	(b"10111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111000100011110101110000101", b"10111111110001010001111010111000"), -- -0.97 + -0.57 = -1.54
	(b"10111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111100110101110000101001000"), -- -0.51 + -0.7 = -1.21
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"10111111011110101110000101001000"), -- -0.54 + -0.44 = -0.98
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"10111110001000111101011100001010"), -- -0.04 + -0.12 = -0.16
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"00111111100011001100110011001101"), -- 0.27 + 0.83 = 1.1
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111100100001010001111010111"), -- 0.23 + 0.9 = 1.13
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110011010111000010100011111", b"10111110111010111000010100011111"), -- -0.23 + -0.23 = -0.46
	(b"10111100101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000111101011100001010010"), -- -0.02 + -0.6 = -0.62
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111011110000101000111101100", b"10111111100110011001100110011010"), -- -0.23 + -0.97 = -1.2

	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000000110011001100110011010"), -- -0.5 + -1.9 = -2.4
	(b"11000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000010101100110011001100110", b"11000000111001110101110000101001"), -- -3.88 + -3.35 = -7.23
	(b"01000000010011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110111100001010001111010111", b"01000000001100010100011110101110"), -- 3.24 + -0.47 = 2.77
	(b"11000000011100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110010101110000101000111101", b"11000000100000001010001111010111"), -- -3.81 + -0.21 = -4.02
	(b"10111111111001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111100010001111010111000011", b"11000000001110000101000111101100"), -- -1.81 + -1.07 = -2.88
	(b"01000000010010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111000000101000111101011100", b"01000000011010101110000101001000"), -- 3.16 + 0.51 = 3.67
	(b"01000000011100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000000011101011100001010010", b"00111111110000111101011100001010"), -- 3.76 + -2.23 = 1.53
	(b"10111111111000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000000110001111010111000011", b"00111111000111101011100001010100"), -- -1.77 + 2.39 = 0.62
	(b"10111111110001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011111110101110000101001", b"11000000101100001111010111000010"), -- -1.54 + -3.99 = -5.53
	(b"11000000011111110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111000011110101110000101001", b"11000000010110111000010100011111"), -- -3.99 + 0.56 = -3.43
	(b"01000000000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"01000000000111110101110000101001"), -- 2.24 + 0.25 = 2.49
	(b"10111111000111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000001001110000101000111101", b"00111111111111111111111111111111"), -- -0.61 + 2.61 = 2
	(b"00111111100111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000000100111101011100001010", b"01000000011000110011001100110011"), -- 1.24 + 2.31 = 3.55
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111110111010111000010100100", b"00111111110010111000010100011111"), -- -0.14 + 1.73 = 1.59
	(b"01000000010100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000011000010100011110101110", b"01000000110110101000111101011100"), -- 3.31 + 3.52 = 6.83
	(b"11000000001101111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010001111010111000010100", b"11000000101111111010111000010100"), -- -2.87 + -3.12 = -5.99
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000101100000000000000000000"), -- 2.8 + 2.7 = 5.5
	(b"10111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111101010001111010111000011", b"10111111111100011110101110000110"), -- -0.57 + -1.32 = -1.89
	(b"01000000010000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111101000111101011100001010", b"00111111110111101011100001010010"), -- 3.02 + -1.28 = 1.74
	(b"11000000000110111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111111011100001010001111011", b"10111111000100011110101110000110"), -- -2.43 + 1.86 = -0.57
	(b"00111111111011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000011000001010001111010111", b"01000000101011000010100011110110"), -- 1.87 + 3.51 = 5.38
	(b"00111111100010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111101011001100110011001101", b"10111110100001010001111010111000"), -- 1.09 + -1.35 = -0.26
	(b"00111111101101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111101010001111010111000010"), -- 1.42 + -0.1 = 1.32
	(b"10111111100010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111110110000101000111101100", b"00111111000110011001100110011010"), -- -1.09 + 1.69 = 0.6
	(b"01000000010100101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111100100001010001111010111", b"01000000100011010111000010100100"), -- 3.29 + 1.13 = 4.42
	(b"00111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110010101110000101000111101", b"00111110101100110011001100110011"), -- 0.14 + 0.21 = 0.35
	(b"10111111101100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000001110101110000101001000", b"11000000100010011001100110011010"), -- -1.38 + -2.92 = -4.3
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000011110101110000101", b"00111110000001010001111010111000"), -- -1.9 + 2.03 = 0.13
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001010001111010111000", b"01000000100111000010100011110110"), -- 2.3 + 2.58 = 4.88
	(b"01000000001100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"00111111111010100011110101110000"), -- 2.78 + -0.95 = 1.83
	(b"00111111100110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111101010100011110101110001", b"10111101111101011100001010010000"), -- 1.21 + -1.33 = -0.12
	(b"01000000011101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111101101011100001010001111", b"01000000101001111010111000010100"), -- 3.82 + 1.42 = 5.24
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111110101000111101011100001", b"00111111100101110000101000111101"), -- -0.48 + 1.66 = 1.18
	(b"10111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111110001110000101000111101100", b"10111100111101011100001010001000"), -- -0.21 + 0.18 = -0.03
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"10111101101000111101011100001000"), -- 0.3 + -0.38 = -0.08
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000011011101011100001010010", b"01000000010111001100110011001101"), -- -0.28 + 3.73 = 3.45
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111111100011110101110000101", b"01000000001010000101000111101100"), -- 0.74 + 1.89 = 2.63
	(b"01000000010010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"01000000010011000010100011110110"), -- 3.15 + 0.04 = 3.19
	(b"11000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"11000000000101011100001010001111"), -- -2.82 + 0.48 = -2.34
	(b"01000000000000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111001001100110011001100110", b"00111111101011100001010001111011"), -- 2.01 + -0.65 = 1.36
	(b"00111111100101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111111110101110000101001000", b"10111111010011001100110011001110"), -- 1.16 + -1.96 = -0.8
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000010000111101011100001010", b"11000000010011100001010001111011"), -- -0.16 + -3.06 = -3.22
	(b"00111111100011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000100011010111000010100100"), -- 1.12 + 3.3 = 4.42
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00111110110001111010111000010101"), -- 0.79 + -0.4 = 0.39
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001010111000010100011111", b"10111111100101011100001010010000"), -- -0.5 + -0.67 = -1.17
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111101111101011100001010001100"), -- -0.52 + 0.4 = -0.12
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010111000010100011110110", b"01000000001101110000101000111110"), -- 2 + 0.86 = 2.86
	(b"10111111101001111010111000010100", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111101001111010111000010100"), -- -1.31 + -0 = -1.31
	(b"10111111111011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111101000000000000000000000", b"11000000010001111010111000010100"), -- -1.87 + -1.25 = -3.12
	(b"00111111111011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000000100011110101110000101", b"10111110110100011110101110000100"), -- 1.87 + -2.28 = -0.41
	(b"11000000011011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111001110000101000111101100", b"11000000010000010100011110101110"), -- -3.74 + 0.72 = -3.02
	(b"10111111110111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111110011100001010001111011", b"10111101111101011100001010010000"), -- -1.73 + 1.61 = -0.12
	(b"11000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"10111111110110011001100110011010"), -- -2.49 + 0.79 = -1.7
	(b"00111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111101111000010100011110101110", b"00111111011100110011001100110011"), -- 0.84 + 0.11 = 0.95
	(b"10111111111010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000000111110101110000101001", b"00111111001001100110011001100110"), -- -1.84 + 2.49 = 0.65
	(b"01000000001101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"01000000010110000101000111101011"), -- 2.86 + 0.52 = 3.38
	(b"01000000000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100000000000000000000", b"10111111100110011001100110011010"), -- 2.05 + -3.25 = -1.2
	(b"10111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111100011110101110000101010"), -- -0.58 + 1.7 = 1.12
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000001101100110011001100110", b"11000000001101110000101000111101"), -- -0.01 + -2.85 = -2.86
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010101011100001010001111", b"11000000011101011100001010001111"), -- -0.5 + -3.34 = -3.84
	(b"11000000010001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010011000010100011110110", b"11000000110010011110101110000101"), -- -3.12 + -3.19 = -6.31
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011100001010001111011", b"00111111010100011110101110000100"), -- -2.9 + 3.72 = 0.82
	(b"10111111110100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111101010001111010111000011", b"11000000001111001100110011001101"), -- -1.63 + -1.32 = -2.95
	(b"00111111111001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111101011001100110011001101", b"01000000010010001111010111000010"), -- 1.79 + 1.35 = 3.14
	(b"10111111100111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000011110111000010100011111", b"11000000101001010001111010111000"), -- -1.23 + -3.93 = -5.16
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"10111101100011110101110000110000"), -- -0.72 + 0.65 = -0.0700001
	(b"11000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111011110000101000111101100", b"11000000100011000111101011100010"), -- -3.42 + -0.97 = -4.39
	(b"11000000000010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000010101111010111000010100", b"00111111100111101011100001010000"), -- -2.13 + 3.37 = 1.24
	(b"11000000001111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000000001011100001010001111", b"11000000101000100011110101110000"), -- -2.98 + -2.09 = -5.07
	(b"01000000010101111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010111110101110000101001", b"10111101111101011100001010100000"), -- 3.37 + -3.49 = -0.12
	(b"11000000010111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001111010111000010100100", b"10111110111110101110000101001000"), -- -3.45 + 2.96 = -0.49
	(b"01000000010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111111110101110000101001000", b"01000000101001111010111000010100"), -- 3.28 + 1.96 = 5.24
	(b"11000000001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"11000000000100111101011100001010"), -- -2.56 + 0.25 = -2.31
	(b"11000000010010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110001010001111010111000", b"11000000100101100001010001111011"), -- -3.15 + -1.54 = -4.69
	(b"01000000011001011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111111010100011110101110001", b"01000000101011010111000010100100"), -- 3.59 + 1.83 = 5.42
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"10111111001010111000010100011110"), -- -1 + 0.33 = -0.67
	(b"11000000001111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111100101011100001010001111", b"11000000100000111000010100011111"), -- -2.94 + -1.17 = -4.11
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111001011100001010001111100"), -- 0.52 + -1.2 = -0.68
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000111010011001100110011010"), -- 3.7 + 3.6 = 7.3
	(b"10111111100000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111100101000111101011100001", b"11000000000010101110000101001000"), -- -1.01 + -1.16 = -2.17
	(b"11000000000000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000000101110000101000111101", b"11000000100011010111000010100100"), -- -2.06 + -2.36 = -4.42
	(b"11000000010101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000000101100110011001100110", b"10111111011111010111000010100100"), -- -3.34 + 2.35 = -0.99
	(b"11000000011100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000011100010100011110101110", b"10111101001000111101011100000000"), -- -3.81 + 3.77 = -0.04
	(b"11000000011100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011101000111101011100001", b"11000000111100100011110101110000"), -- -3.75 + -3.82 = -7.57
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000011101010001111010111000", b"11000000010000110011001100110011"), -- 0.78 + -3.83 = -3.05
	(b"10111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"10111110011000010100011110101110"), -- -0.44 + 0.22 = -0.22
	(b"11000000000010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110101000111101011100001010", b"11000000000111100001010001111011"), -- -2.15 + -0.32 = -2.47
	(b"00111111101101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"00111110110111000010100011110100"), -- 1.42 + -0.99 = 0.43
	(b"10111111111001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000011001111010111000010100", b"11000000101011011100001010001111"), -- -1.81 + -3.62 = -5.43
	(b"01000000000111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000010111000010100011110110", b"10111111011101011100001010010000"), -- 2.48 + -3.44 = -0.96
	(b"11000000001001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000011010100011110101110001", b"11000000110010001010001111010111"), -- -2.61 + -3.66 = -6.27
	(b"11000000010010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111111101110000101000111101", b"11000000101000100011110101110001"), -- -3.14 + -1.93 = -5.07
	(b"10111110001011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000010010101110000101001000", b"11000000010101011100001010010000"), -- -0.17 + -3.17 = -3.34
	(b"01000000010001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000011110101110000101001000", b"10111111010011110101110000101100"), -- 3.11 + -3.92 = -0.81
	(b"10111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111110101011100001010001111", b"00111111011010001111010111000010"), -- -0.76 + 1.67 = 0.91
	(b"00111111100010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000010001111010111000010100", b"11000000000000011110101110000100"), -- 1.09 + -3.12 = -2.03
	(b"01000000011000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000011010001111010111000011", b"01000000111001100110011001100110"), -- 3.56 + 3.64 = 7.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000101100110011001100110", b"01000000000101100110011001100110"), -- -0 + 2.35 = 2.35
	(b"10111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000010110100011110101110001", b"01000000010001000111101011100010"), -- -0.34 + 3.41 = 3.07
	(b"11000000001000011110101110000101", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"11000000000111110101110000101001"), -- -2.53 + 0.04 = -2.49
	(b"10111111101111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000010111010111000010100100", b"00111111111111010111000010100100"), -- -1.48 + 3.46 = 1.98
	(b"10111111110111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000000111100001010001111011", b"11000000100001100001010001111011"), -- -1.72 + -2.47 = -4.19
	(b"01000000011011010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000011111000010100011110110", b"10111110011010111000010100100000"), -- 3.71 + -3.94 = -0.23
	(b"11000000000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001110000101000111101100", b"00111111000001111010111000011000"), -- -2.35 + 2.88 = 0.53
	(b"11000000001001110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000010001011100001010001111", b"00111110111101011100001010010000"), -- -2.61 + 3.09 = 0.48
	(b"00111111110100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111111011100001010001111011", b"10111110011010111000010100100000"), -- 1.63 + -1.86 = -0.23
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000001111110101110000101001", b"11000000001011001100110011001101"), -- 0.29 + -2.99 = -2.7
	(b"11000000011111110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111100010001111010111000011", b"11000000001110101110000101001000"), -- -3.99 + 1.07 = -2.92
	(b"00111111111101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111100011100001010001111011", b"00111111010011001100110011001100"), -- 1.91 + -1.11 = 0.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001110000101000111101", b"00111111111001111010111000010100"), -- -0.3 + 2.11 = 1.81
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111111100011110101110000101", b"00111111100010001111010111000010"), -- -0.82 + 1.89 = 1.07
	(b"00111111111110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"01000000000010111000010100011111"), -- 1.94 + 0.24 = 2.18
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111110100010100011110101110001", b"00111110000001010001111010111001"), -- -0.14 + 0.27 = 0.13
	(b"01000000000001011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000001100011110101110000101", b"01000000100110111101011100001010"), -- 2.09 + 2.78 = 4.87
	(b"00111111101010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111111011110101110000101001", b"10111111000010100011110101110000"), -- 1.33 + -1.87 = -0.54
	(b"01000000011010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000000101111010111000010100", b"01000000110000001111010111000010"), -- 3.66 + 2.37 = 6.03
	(b"01000000001000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001011100001010001111", b"01000000101101000111101011100001"), -- 2.55 + 3.09 = 5.64
	(b"01000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000011011110101110000101001", b"01000000110110000000000000000000"), -- 3.01 + 3.74 = 6.75
	(b"11000000001111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000110011001100110011", b"11000000110100000000000000000000"), -- -2.95 + -3.55 = -6.5
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010010001111010111000011", b"11000000011101010001111010111001"), -- -0.69 + -3.14 = -3.83
	(b"00111111111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000110011001100110011", b"10111111001100110011001100110010"), -- 1.85 + -2.55 = -0.7
	(b"00111111111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011101010001111010111000", b"10111111111100001010001111010110"), -- 1.95 + -3.83 = -1.88
	(b"10111111110000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111100010111000010100011111", b"10111110111000010100011110101100"), -- -1.53 + 1.09 = -0.44
	(b"11000000000001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000000100101000111101011100", b"00111110010101110000101001000000"), -- -2.08 + 2.29 = 0.21
	(b"11000000001110100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111111101000111101011100001", b"11000000100110100011110101110001"), -- -2.91 + -1.91 = -4.82
	(b"00111111110101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000000011000010100011110110", b"01000000011101110000101000111110"), -- 1.67 + 2.19 = 3.86
	(b"11000000010111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100101110000101000111101", b"11000000100101000010100011110110"), -- -3.45 + -1.18 = -4.63
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011010001111010111000011", b"01000000110010101110000101001000"), -- 2.7 + 3.64 = 6.34
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000010010111000010100011111", b"11000000000110001111010111000011"), -- 0.79 + -3.18 = -2.39
	(b"01000000010011000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"01000000000101011100001010010000"), -- 3.19 + -0.85 = 2.34
	(b"10111111100010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"10111111010100011110101110000110"), -- -1.07 + 0.25 = -0.82
	(b"11000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"11000000010011001100110011001101"), -- -2.42 + -0.78 = -3.2
	(b"00111111110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000010000101000111101100", b"10111110111101011100001010010100"), -- 1.65 + -2.13 = -0.48
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101011100001010001111011", b"00111111101011100001010001111011"), -- -0 + 1.36 = 1.36
	(b"01000000000011000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111111101011100001010001111", b"01000000100000111000010100011111"), -- 2.19 + 1.92 = 4.11
	(b"01000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111111000111101011100001010", b"01000000101001100110011001100110"), -- 3.42 + 1.78 = 5.2
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111111101011100001010001111", b"10111111110001010001111010111000"), -- 0.38 + -1.92 = -1.54
	(b"00111111101101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111110111000010100011110110"), -- 1.42 + 0.3 = 1.72
	(b"11000000011111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011111010111000010100100", b"00111100001000111101011100000000"), -- -3.95 + 3.96 = 0.00999999
	(b"00111111100000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111010000101000111101011100", b"00111110100010100011110101110000"), -- 1.03 + -0.76 = 0.27
	(b"01000000010101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000011001000111101011100001", b"01000000110111011100001010001111"), -- 3.36 + 3.57 = 6.93
	(b"01000000001000011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101000001111010111000010"), -- 2.53 + 2.5 = 5.03
	(b"01000000001000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001110000101000111101", b"01000000110001010001111010111000"), -- 2.55 + 3.61 = 6.16
	(b"11000000010011000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111110010111000010100011111", b"10111111110011001100110011001101"), -- -3.19 + 1.59 = -1.6
	(b"00111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000011011110101110000101001", b"11000000010101111010111000010100"), -- 0.37 + -3.74 = -3.37
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000001011101011100001010010"), -- -0.87 + 3.6 = 2.73
	(b"01000000001101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011011110101110000101001", b"01000000110100101110000101001000"), -- 2.85 + 3.74 = 6.59
	(b"10111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111111101110000101000111101", b"00111111101011001100110011001100"), -- -0.58 + 1.93 = 1.35
	(b"11000000010010101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000011010101110000101001000", b"11000000110110101110000101001000"), -- -3.17 + -3.67 = -6.84
	(b"00111110000001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011100101000111101011100", b"11000000011010100011110101110000"), -- 0.13 + -3.79 = -3.66
	(b"01000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111111100001010001111010111", b"00111111110001010001111010111001"), -- 3.42 + -1.88 = 1.54
	(b"10111111101000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111101101110000101000111101", b"11000000001011001100110011001100"), -- -1.27 + -1.43 = -2.7
	(b"11000000010011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111110100001010001111010111", b"11000000100110110011001100110011"), -- -3.22 + -1.63 = -4.85
	(b"11000000001011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000000011101011100001010010", b"11000000100111100110011001100110"), -- -2.72 + -2.23 = -4.95
	(b"11000000011110100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000001010011001100110011010", b"10111111101000010100011110101110"), -- -3.91 + 2.65 = -1.26
	(b"11000000001010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111110011110101110000101001", b"10111111100000101000111101011101"), -- -2.64 + 1.62 = -1.02
	(b"10111111111110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"10111111110001111010111000010101"), -- -1.95 + 0.39 = -1.56
	(b"00111111010000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000001110111000010100011111", b"01000000011011000010100011110110"), -- 0.76 + 2.93 = 3.69
	(b"10111111110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000101010110011001100110011"), -- -1.65 + -3.7 = -5.35
	(b"10111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111100010001111010111000011", b"10111111110110011001100110011010"), -- -0.63 + -1.07 = -1.7
	(b"11000000000101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"10111111110110000101000111101011"), -- -2.34 + 0.65 = -1.69
	(b"10111111101010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000011110000101000111101100", b"11000000101001110000101000111110"), -- -1.34 + -3.88 = -5.22
	(b"01000000001111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000000111101011100001010010", b"01000000101011110000101000111110"), -- 2.99 + 2.48 = 5.47
	(b"00111111101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100111100110011001100110"), -- 1.45 + 3.5 = 4.95
	(b"11000000001001000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000011001000111101011100001"), -- -2.57 + -1 = -3.57
	(b"11000000011110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"11000000010111010111000010100100"), -- -3.92 + 0.46 = -3.46
	(b"10111111110001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111111101110000101000111101", b"00111110110001111010111000010100"), -- -1.54 + 1.93 = 0.39
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"11000000001000000000000000000000"), -- -2.4 + -0.1 = -2.5
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000101100110011001100110", b"11000000101110110011001100110011"), -- -3.5 + -2.35 = -5.85
	(b"10111111110110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000010011101011100001010010", b"11000000100111010111000010100100"), -- -1.69 + -3.23 = -4.92
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001111100001010001111011", b"01000000011101110000101000111110"), -- 0.89 + 2.97 = 3.86
	(b"01000000010100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000010001110000101000111101", b"01000000110010111101011100001010"), -- 3.26 + 3.11 = 6.37
	(b"00111111100101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111100011100001010001111011", b"01000000000100101000111101011100"), -- 1.18 + 1.11 = 2.29
	(b"01000000001110001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000011110000101000111101100", b"01000000110110001010001111011000"), -- 2.89 + 3.88 = 6.77
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011010011001100110011010"), -- 0.05 + -3.7 = -3.65
	(b"10111111101101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000010010101110000101001000", b"00111111110111101011100001010011"), -- -1.43 + 3.17 = 1.74
	(b"11000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000010101111010111000010100", b"11000000110010011001100110011010"), -- -2.93 + -3.37 = -6.3
	(b"11000000010101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000010011101011100001010010", b"11000000110100100011110101110000"), -- -3.34 + -3.23 = -6.57
	(b"10111110111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101001010001111010111000", b"10111111110111101011100001010010"), -- -0.45 + -1.29 = -1.74
	(b"00111111100111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000010100011110101110000101", b"01000000100100000000000000000000"), -- 1.22 + 3.28 = 4.5
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000101000111101011100", b"10111110111010111000010100100000"), -- -3.5 + 3.04 = -0.46
	(b"00111111110100011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000011111100001010001111011", b"01000000101100111000010100011111"), -- 1.64 + 3.97 = 5.61
	(b"01000000001010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110100110011001100110011", b"00111111100000000000000000000001"), -- 2.65 + -1.65 = 1
	(b"00111111110100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111110100110011001100110011", b"10111100101000111101011100000000"), -- 1.63 + -1.65 = -0.02
	(b"10111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111101111010111000010100100", b"00111111101101011100001010010000"), -- -0.06 + 1.48 = 1.42
	(b"01000000010011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000011000110011001100110011", b"10111110101010001111010111000000"), -- 3.22 + -3.55 = -0.33
	(b"10111111101111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000000001011100001010001111", b"11000000011001010001111010111000"), -- -1.49 + -2.09 = -3.58
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111111100011110101110000101", b"10111111110000111101011100001010"), -- 0.36 + -1.89 = -1.53
	(b"10111111111011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000101000111101011100001", b"10111111101000101000111101011100"), -- -1.85 + 0.58 = -1.27
	(b"10111111111110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000011010111000010100011111", b"00111111110111101011100001010010"), -- -1.94 + 3.68 = 1.74
	(b"11000000000110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000010101010001111010111000", b"00111111011100110011001100110000"), -- -2.38 + 3.33 = 0.95
	(b"00111111110111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000001101000111101011100001", b"01000000100100011110101110000101"), -- 1.74 + 2.82 = 4.56
	(b"10111111110111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000000110000101000111101100", b"11000000100000110011001100110100"), -- -1.72 + -2.38 = -4.1
	(b"10111111100110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111110101110000101000111101", b"11000000001110001111010111000010"), -- -1.21 + -1.68 = -2.89
	(b"10111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"10111110110100011110101110000100"), -- -0.58 + 0.17 = -0.41
	(b"00111111110110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111111000101110000101000111100"), -- 1.71 + -2.3 = -0.59
	(b"10111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000000001110000101000111101", b"11000000001101100110011001100110"), -- -0.74 + -2.11 = -2.85
	(b"00111111101110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"00111111000011110101110000101010"), -- 1.45 + -0.89 = 0.56
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"10111110010101110000101000111101"), -- -0.16 + -0.05 = -0.21
	(b"10111111100001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000011011110101110000101001", b"01000000001011001100110011001101"), -- -1.04 + 3.74 = 2.7
	(b"10111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"10111111010000101000111101011100"), -- -0.73 + -0.03 = -0.76
	(b"01000000000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110111000010100011111", b"01000000101011110101110000101001"), -- 2.05 + 3.43 = 5.48
	(b"11000000001100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111110101011100001010001111", b"11000000100011100110011001100110"), -- -2.78 + -1.67 = -4.45
	(b"10111111100001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011000110011001100110011", b"11000000100100101110000101001000"), -- -1.04 + -3.55 = -4.59
	(b"11000000001000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111001101011100001010001111", b"10111111111010100011110101110000"), -- -2.54 + 0.71 = -1.83
	(b"01000000011000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"01000000001011101011100001010010"), -- 3.51 + -0.78 = 2.73
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011000010100011110110"), -- -0.01 + 2.2 = 2.19
	(b"00111111111111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111101010111000010100011111", b"01000000010100111101011100001010"), -- 1.97 + 1.34 = 3.31
	(b"10111111101010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000010001000111101011100001", b"11000000100011000111101011100001"), -- -1.32 + -3.07 = -4.39
	(b"01000000011000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000011011000010100011110110", b"01000000111001110101110000101001"), -- 3.54 + 3.69 = 7.23
	(b"01000000010001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000010100111101011100001010", b"10111110010011001100110011010000"), -- 3.11 + -3.31 = -0.2
	(b"00111111000011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000010101010001111010111000", b"01000000011110001111010111000010"), -- 0.56 + 3.33 = 3.89
	(b"11000000000001000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111100010111000010100011111", b"11000000010010100011110101110000"), -- -2.07 + -1.09 = -3.16
	(b"10111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000011101100110011001100110", b"01000000010001111010111000010100"), -- -0.73 + 3.85 = 3.12
	(b"00111111110111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000000101000111101011100001", b"10111111000101000111101011100000"), -- 1.74 + -2.32 = -0.58
	(b"01000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000000100010100011110101110"), -- 2.97 + -0.7 = 2.27
	(b"11000000011101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111110010100011110101110001", b"11000000000100011110101110000100"), -- -3.86 + 1.58 = -2.28
	(b"11000000000100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101010001111010111000011", b"11000000011001000111101011100010"), -- -2.25 + -1.32 = -3.57
	(b"10111111111110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000001110100011110101110001", b"00111111011100110011001100110100"), -- -1.96 + 2.91 = 0.95
	(b"11000000001100101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111101100001010001111010111", b"11000000100001010111000010100100"), -- -2.79 + -1.38 = -4.17
	(b"00111111101100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000010101010001111010111000", b"01000000100101101011100001010010"), -- 1.38 + 3.33 = 4.71
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110101000111101011100001010", b"01000000100000001010001111010111"), -- 3.7 + 0.32 = 4.02
	(b"00111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000010001010001111010111000", b"01000000100000011001100110011010"), -- 0.97 + 3.08 = 4.05
	(b"11000000001111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001111010111000010100", b"11000000100010000101000111101100"), -- -2.95 + -1.31 = -4.26
	(b"10111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111001101011100001010001111", b"10111111100111010111000010100100"), -- -0.52 + -0.71 = -1.23
	(b"00111111101111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"00111111001001100110011001100111"), -- 1.48 + -0.83 = 0.65
	(b"11000000000110100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111101001010001111010111000", b"11000000011011001100110011001101"), -- -2.41 + -1.29 = -3.7
	(b"01000000011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111101000101000111101011100", b"01000000100110010100011110101110"), -- 3.52 + 1.27 = 4.79
	(b"11000000011001000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111010001111010111000010100", b"11000000001100101000111101011100"), -- -3.57 + 0.78 = -2.79
	(b"11000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000010110100011110101110000"), -- -2.81 + -0.6 = -3.41
	(b"11000000000101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111100000101000111101011100", b"10111111101001100110011001100110"), -- -2.32 + 1.02 = -1.3
	(b"10111111111101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000001110100011110101110001", b"11000000100110100011110101110001"), -- -1.91 + -2.91 = -4.82
	(b"01000000011010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"00111111100001111010111000010110"), -- 3.66 + -2.6 = 1.06
	(b"01000000011100010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000010010000101000111101100", b"01000000110111001100110011001101"), -- 3.77 + 3.13 = 6.9
	(b"10111111100100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110110101110000101000111101", b"10111111001101011100001010010000"), -- -1.13 + 0.42 = -0.71
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110100011110101110001", b"11000000110011010001111010111000"), -- -3.5 + -2.91 = -6.41
	(b"11000000010100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000110010001111010111000010"), -- -3.28 + -3 = -6.28
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000000000110011001100110011", b"00111111111000101000111101011100"), -- -0.28 + 2.05 = 1.77
	(b"10111111111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111111110000101000111101100", b"00111100101000111101011101000000"), -- -1.92 + 1.94 = 0.0200001
	(b"11000000001111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010111010111000010100100", b"11000000110011010001111010111000"), -- -2.95 + -3.46 = -6.41
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000011000010100011110110", b"00111110100101000111101011100100"), -- -1.9 + 2.19 = 0.29
	(b"10111110110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111111011110101110000101001", b"00111111101110101110000101001000"), -- -0.41 + 1.87 = 1.46
	(b"10111111100110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000011100010100011110101110", b"01000000001000111101011100001010"), -- -1.21 + 3.77 = 2.56
	(b"11000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000000011010111000010100100", b"10111110100011110101110000101000"), -- -2.49 + 2.21 = -0.28
	(b"00111111100101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000011001010001111010111000"), -- 1.18 + 2.4 = 3.58
	(b"10111111011110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000001101111010111000010100", b"00111111111100011110101110000100"), -- -0.98 + 2.87 = 1.89
	(b"00111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111110111101011100001010010", b"01000000000110111000010100011111"), -- 0.69 + 1.74 = 2.43
	(b"01000000011010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000101000111101011100001", b"01000000101111110000101000111110"), -- 3.65 + 2.32 = 5.97
	(b"10111111110000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111111111010111000010100100", b"11000000011000000000000000000000"), -- -1.52 + -1.98 = -3.5
	(b"10111111110010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000011011010111000010100100", b"01000000000010001111010111000010"), -- -1.57 + 3.71 = 2.14
	(b"10111111111000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000100001010111000010100100"), -- -1.77 + -2.4 = -4.17
	(b"01000000000100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101110000101000111101100", b"01000000011011000010100011110110"), -- 2.25 + 1.44 = 3.69
	(b"10111111111011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000001101010001111010111000", b"11000000100101100110011001100110"), -- -1.87 + -2.83 = -4.7
	(b"10111111100000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000010011110101110000101001", b"01000000000011010111000010100100"), -- -1.03 + 3.24 = 2.21
	(b"00111110111100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111110111010111000010100011111", b"00111100001000111101011100000000"), -- 0.47 + -0.46 = 0.00999999
	(b"11000000010110001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000010101100110011001100110", b"11000000110101111010111000010100"), -- -3.39 + -3.35 = -6.74
	(b"11000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111010000000000000000000000", b"11000000010011110101110000101001"), -- -2.49 + -0.75 = -3.24
	(b"11000000011100101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000001000010100011110101110", b"10111111101000101000111101011100"), -- -3.79 + 2.52 = -1.27
	(b"01000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"01000000010111010111000010100100"), -- 3.01 + 0.45 = 3.46
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"11000000011100111101011100001010"), -- -3.8 + -0.01 = -3.81
	(b"01000000010001110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111111000010100011110101110", b"00111111101011001100110011001100"), -- 3.11 + -1.76 = 1.35
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"00111111100000010100011110101110"), -- 0.34 + 0.67 = 1.01
	(b"10111111101010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111111101000111101011100010"), -- -1.32 + -0.59 = -1.91
	(b"10111111101001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010111010111000010100100", b"11000000100110001010001111010111"), -- -1.31 + -3.46 = -4.77
	(b"11000000000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111100100011110101110000101", b"11000000011001111010111000010100"), -- -2.48 + -1.14 = -3.62
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110011010111000010100011111", b"10111111110101011100001010001111"), -- -1.9 + 0.23 = -1.67
	(b"11000000011001011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111101011001100110011001101", b"11000000100111100001010001111011"), -- -3.59 + -1.35 = -4.94
	(b"01000000011000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000100100111000010100011111"), -- 3.51 + 1.1 = 4.61
	(b"01000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000000110111000010100011111", b"01000000101010000000000000000000"), -- 2.82 + 2.43 = 5.25
	(b"11000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000000111100001010001111011", b"11000000110010110011001100110100"), -- -3.88 + -2.47 = -6.35
	(b"11000000010011010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111110111010111000010100100", b"11000000100111100001010001111011"), -- -3.21 + -1.73 = -4.94
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001010001111010111000", b"00111111011110101110000101001000"), -- -2.6 + 3.58 = 0.98
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000010100011110101110", b"01000000000011100001010001111011"), -- -0.3 + 2.52 = 2.22
	(b"11000000011000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111101101000111101011100001010", b"11000000010111101011100001010010"), -- -3.56 + 0.08 = -3.48
	(b"01000000010011101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111001110101110000101001000"), -- 3.23 + -2.5 = 0.73
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010111000010100011110110", b"10111111101000010100011110101110"), -- -0.4 + -0.86 = -1.26
	(b"11000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000010100001010001111010111", b"11000000110001100001010001111011"), -- -2.93 + -3.26 = -6.19
	(b"10111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000011011110101110000101001", b"01000000011010011001100110011010"), -- -0.09 + 3.74 = 3.65
	(b"01000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111111000101110000101000111100"), -- 2.51 + -3.1 = -0.59
	(b"11000000000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"11000000010100110011001100110011"), -- -2.48 + -0.82 = -3.3
	(b"10111111110101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111111111010111000010100100", b"00111110100111101011100001010100"), -- -1.67 + 1.98 = 0.31
	(b"00111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010010101110000101001000"), -- 0.03 + -3.2 = -3.17
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001110000101000111101100", b"00111111111111101011100001010011"), -- -0.89 + 2.88 = 1.99
	(b"00111111111111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111100010111000010100011111", b"00111111011001100110011001100110"), -- 1.99 + -1.09 = 0.9
	(b"01000000010111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111100011100001010001111011", b"01000000000101100110011001100110"), -- 3.46 + -1.11 = 2.35
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000000111110101110000101001", b"11000000001111101011100001010010"), -- -0.49 + -2.49 = -2.98
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"11000000000000110011001100110011"), -- -2.3 + 0.25 = -2.05
	(b"00111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111111111000010100011110110", b"10111111101001111010111000010100"), -- 0.66 + -1.97 = -1.31
	(b"11000000011001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111000101110000101000111101", b"11000000010000011110101110000101"), -- -3.62 + 0.59 = -3.03
	(b"10111111101101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000010010000101000111101100", b"00111111110110101110000101001001"), -- -1.42 + 3.13 = 1.71
	(b"10111100111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111110011100001010001111011", b"10111111110100011110101110000101"), -- -0.03 + -1.61 = -1.64
	(b"10111111101011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"10111111100101110000101000111110"), -- -1.35 + 0.17 = -1.18
	(b"01000000010110100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000000000110011001100110011", b"01000000101011101011100001010010"), -- 3.41 + 2.05 = 5.46
	(b"01000000000101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000010111110101110000101001", b"10111111100100001010001111011000"), -- 2.36 + -3.49 = -1.13
	(b"11000000011000011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000001101100110011001100110", b"11000000110011000010100011110110"), -- -3.53 + -2.85 = -6.38
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000000001010001111010111000", b"00111111100111101011100001010010"), -- -0.84 + 2.08 = 1.24
	(b"01000000001100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"01000000001011110101110000101001"), -- 2.78 + -0.04 = 2.74
	(b"10111111111010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110111001100110011001100110", b"10111111101011110101110000101010"), -- -1.82 + 0.45 = -1.37
	(b"11000000001010101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000011010111000010100011111", b"11000000110010110011001100110100"), -- -2.67 + -3.68 = -6.35
	(b"11000000011110001111010111000011", b"00000000000000000000000000000000"),
	(b"00111110011000010100011110101110", b"11000000011010101110000101001000"), -- -3.89 + 0.22 = -3.67
	(b"11000000010101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110101010001111010111000011", b"11000000001111110101110000101001"), -- -3.32 + 0.33 = -2.99
	(b"10111111100100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010110111000010100011111", b"11000000100100011110101110000101"), -- -1.13 + -3.43 = -4.56
	(b"10111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000001101111010111000010100", b"11000000010100110011001100110011"), -- -0.43 + -2.87 = -3.3
	(b"11000000011000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010000000000000000000000", b"11000000001100110011001100110011"), -- -3.55 + 0.75 = -2.8
	(b"01000000000001110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111110000010100011110101101"), -- 2.11 + -0.6 = 1.51
	(b"11000000011100011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111111000111101011100001010"), -- -3.78 + 2 = -1.78
	(b"01000000010111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000011001111010111000010100", b"10111110001110000101000111100000"), -- 3.44 + -3.62 = -0.18
	(b"00111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111111001111010111000010100", b"01000000000001100110011001100110"), -- 0.29 + 1.81 = 2.1
	(b"01000000010010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"01000000001110001111010111000011"), -- 3.15 + -0.26 = 2.89
	(b"00111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000000100101000111101011100", b"10111111111011001100110011001100"), -- 0.44 + -2.29 = -1.85
	(b"01000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111110100101000111101011100000"), -- 2.51 + -2.8 = -0.29
	(b"10111111101001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111101111000010100011110101110", b"10111111100110011001100110011001"), -- -1.31 + 0.11 = -1.2
	(b"01000000011111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011100001010001111011", b"01000000001101011100001010010000"), -- 3.95 + -1.11 = 2.84
	(b"10111111101001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111101010011001100110011001101", b"10111111101000010100011110101110"), -- -1.31 + 0.05 = -1.26
	(b"11000000011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110000011110101110000101001", b"11000000011010100011110101110001"), -- -3.52 + -0.14 = -3.66
	(b"11000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000001111001100110011001101", b"11000000110100001111010111000010"), -- -3.58 + -2.95 = -6.53
	(b"11000000010010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000010011110101110000101001", b"11000000110011010111000010100100"), -- -3.18 + -3.24 = -6.42
	(b"10111111110110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000010110101110000101001000", b"11000000101001000010100011110110"), -- -1.71 + -3.42 = -5.13
	(b"11000000011001000111101011100001", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"11000000011001110000101000111101"), -- -3.57 + -0.04 = -3.61
	(b"11000000001001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000001110000101000111101100", b"00111110100110011001100110100000"), -- -2.58 + 2.88 = 0.3
	(b"11000000010110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000001011100001010001111011", b"11000000110001001100110011001101"), -- -3.43 + -2.72 = -6.15
	(b"00111111110101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111101110000101000111101100", b"00111110011101011100001010001000"), -- 1.68 + -1.44 = 0.24
	(b"10111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000000000111101011100001010", b"11000000010000110011001100110011"), -- -0.99 + -2.06 = -3.05
	(b"01000000000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011101010001111010111000", b"10111111101111010111000010100100"), -- 2.35 + -3.83 = -1.48
	(b"11000000000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111101100011110101110000101", b"10111111010110011001100110011010"), -- -2.24 + 1.39 = -0.85
	(b"01000000010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111110111101011100001010010", b"00111111110011110101110000101000"), -- 3.36 + -1.74 = 1.62
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011010111000010100100", b"00111111010010100011110101110000"), -- 3 + -2.21 = 0.79
	(b"00111111100100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000011011100001010001111011", b"11000000001001011100001010010000"), -- 1.13 + -3.72 = -2.59
	(b"00111111101010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000011000011110101110000110"), -- 1.33 + 2.2 = 3.53
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000011101110000101000111101", b"11000000100000000000000000000000"), -- -0.14 + -3.86 = -4
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000011010111000010100011111", b"01000000011110001111010111000011"), -- 0.21 + 3.68 = 3.89
	(b"00111111100110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000001111100001010001111011", b"01000000100001010001111010111000"), -- 1.19 + 2.97 = 4.16
	(b"00111111101110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"00111111111101000111101011100010"), -- 1.45 + 0.46 = 1.91
	(b"01000000001101010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000001010001111010111000011", b"01000000101011110000101000111110"), -- 2.83 + 2.64 = 5.47
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011010111000010100100", b"01000000100011010001111010111000"), -- 2.2 + 2.21 = 4.41
	(b"10111111111110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100000010100011110101110", b"10111111011100001010001111011000"), -- -1.95 + 1.01 = -0.94
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010110011001100110011010", b"11000000010111001100110011001100"), -- -2.6 + -0.85 = -3.45
	(b"00111111000101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000011110100011110101110001", b"01000000100011111010111000010101"), -- 0.58 + 3.91 = 4.49
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"10111111001010001111010111000010"), -- -0.25 + -0.41 = -0.66
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000011010000101000111101100"), -- 0.23 + 3.4 = 3.63
	(b"01000000001101010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000011110100011110101110001", b"01000000110101111010111000010100"), -- 2.83 + 3.91 = 6.74
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000010100000000000000000000", b"11000000011011101011100001010010"), -- -0.48 + -3.25 = -3.73
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011101100110011001100110", b"11000000111100011001100110011010"), -- -3.7 + -3.85 = -7.55
	(b"10111111111000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111111011110101110000101000111"), -- -1.78 + 0.8 = -0.98
	(b"10111111100111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"10111111011111010111000010100100"), -- -1.24 + 0.25 = -0.99
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111001110000101000111101100", b"10111111110001111010111000010100"), -- -0.84 + -0.72 = -1.56
	(b"10111111101000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111010001111010111000011", b"11000000010001000111101011100010"), -- -1.25 + -1.82 = -3.07
	(b"00111111101011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111110000101000111101100", b"01000000010100101000111101011100"), -- 1.35 + 1.94 = 3.29
	(b"11000000010100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"11000000011001011100001010001111"), -- -3.26 + -0.33 = -3.59
	(b"11000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110110000101000111101011100", b"11000000000000101000111101011100"), -- -2.42 + 0.38 = -2.04
	(b"10111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000001101000111101011100001", b"11000000010010100011110101110000"), -- -0.34 + -2.82 = -3.16
	(b"10111111101101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"00111111000101110000101000111110"), -- -1.41 + 2 = 0.59
	(b"00111110101010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111100001010001111010111000", b"10111111001101011100001010001110"), -- 0.33 + -1.04 = -0.71
	(b"01000000000111100001010001111011", b"00000000000000000000000000000000"),
	(b"00111101111101011100001010001111", b"01000000001001011100001010001111"), -- 2.47 + 0.12 = 2.59
	(b"01000000000100101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111111001111010111000010100", b"01000000100000110011001100110011"), -- 2.29 + 1.81 = 4.1
	(b"00111111110100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000001101100110011001100110", b"01000000100011110101110000101001"), -- 1.63 + 2.85 = 4.48
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000000010001111010111000011", b"00111111110011100001010001111100"), -- -0.53 + 2.14 = 1.61
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000000010101110000101001000", b"11000000010000101000111101011100"), -- -0.87 + -2.17 = -3.04
	(b"11000000001010101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000011111101011100001010010", b"11000000110101001100110011001101"), -- -2.67 + -3.98 = -6.65
	(b"11000000000001110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000000101010001111010111000", b"00111110011000010100011110110000"), -- -2.11 + 2.33 = 0.22
	(b"01000000010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"01000000010100111101011100001010"), -- 3.24 + 0.07 = 3.31
	(b"10111111110010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000010101111010111000010100", b"11000000100111100110011001100110"), -- -1.58 + -3.37 = -4.95
	(b"11000000000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000101000111101011100001", b"11000000100100100011110101110000"), -- -2.25 + -2.32 = -4.57
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000010000110011001100110011", b"11000000000111010111000010100100"), -- 0.59 + -3.05 = -2.46
	(b"10111111101010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000010011000010100011110110", b"00111111111011001100110011001101"), -- -1.34 + 3.19 = 1.85
	(b"11000000001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"11000000000110100011110101110001"), -- -2.88 + 0.47 = -2.41
	(b"11000000011010000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111100110101110000101001000", b"11000000000110101110000101001000"), -- -3.63 + 1.21 = -2.42
	(b"11000000001011010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000011111101011100001010010", b"11000000110101100001010001111011"), -- -2.71 + -3.98 = -6.69
	(b"10111111100101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111111011110101110000101001", b"00111111001101011100001010010000"), -- -1.16 + 1.87 = 0.71
	(b"11000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000011010000101000111101100", b"10111110101100110011001100110000"), -- -3.98 + 3.63 = -0.35
	(b"10111111100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111101000000000000000000000"), -- -1.05 + 2.3 = 1.25
	(b"10111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"00111101101000111101011100001000"), -- -0.54 + 0.62 = 0.08
	(b"11000000000011000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"11000000000101100110011001100111"), -- -2.19 + -0.16 = -2.35
	(b"11000000011101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001111010111000010100", b"10111111001110101110000101001000"), -- -3.85 + 3.12 = -0.73
	(b"00111111110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010010100011110101110001", b"01000000100101101011100001010010"), -- 1.55 + 3.16 = 4.71
	(b"00111110010101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111000100011110101110000101", b"00111111010001111010111000010100"), -- 0.21 + 0.57 = 0.78
	(b"11000000010110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000011010011001100110011010", b"00111110100010100011110101110000"), -- -3.38 + 3.65 = 0.27
	(b"10111111110111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000001101000111101011100001", b"00111111100011001100110011001100"), -- -1.72 + 2.82 = 1.1
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"10111111100000000000000000000000"), -- -3.7 + 2.7 = -1
	(b"11000000010101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001011100001010001111", b"10111111101000010100011110101110"), -- -3.35 + 2.09 = -1.26
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000001000110011001100110011", b"11000000010101110000101000111101"), -- -0.81 + -2.55 = -3.36
	(b"11000000001110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000010011010111000010100100", b"00111110101010001111010111000000"), -- -2.88 + 3.21 = 0.33
	(b"10111111101010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111011110101110000101000110"), -- -1.32 + 2.3 = 0.98
	(b"10111111101100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111110001100110011001100110", b"11000000001111000010100011110110"), -- -1.39 + -1.55 = -2.94
	(b"00111111110101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110010000101000111101011100", b"00111111101111010111000010100100"), -- 1.67 + -0.19 = 1.48
	(b"10111111111100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111101101011100001010001111"), -- -1.88 + 3.3 = 1.42
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000000011110101110000101", b"00111111110101011100001010001111"), -- -0.36 + 2.03 = 1.67
	(b"10111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111111000111101011100001010", b"11000000000110100011110101110000"), -- -0.63 + -1.78 = -2.41
	(b"01000000011000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000111110101110000101001", b"00111111100001111010111000010100"), -- 3.55 + -2.49 = 1.06
	(b"10111111101010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111100010001111010111000011", b"11000000000110011001100110011010"), -- -1.33 + -1.07 = -2.4
	(b"01000000011100101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111100000101000111101011100", b"01000000001100010100011110101110"), -- 3.79 + -1.02 = 2.77
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111100101000111101011100001"), -- -0.96 + -0.2 = -1.16
	(b"00111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000001101111010111000010100", b"01000000010000001010001111010111"), -- 0.14 + 2.87 = 3.01
	(b"10111111101111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000000101100110011001100110", b"00111111011000010100011110101100"), -- -1.47 + 2.35 = 0.88
	(b"10111111101010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000001010011001100110011010", b"11000000011111100001010001111100"), -- -1.32 + -2.65 = -3.97
	(b"11000000000001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000001111101011100001010010", b"11000000101000110011001100110011"), -- -2.12 + -2.98 = -5.1
	(b"00111111111010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"00111111110110011001100110011010"), -- 1.82 + -0.12 = 1.7
	(b"01000000010000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101010100011110101110001", b"00111111110111000010100011110101"), -- 3.05 + -1.33 = 1.72
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110111101011100001010001111", b"11000000010001111010111000010100"), -- -3.6 + 0.48 = -3.12
	(b"10111111000100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000010101111010111000010100"), -- -0.57 + -2.8 = -3.37
	(b"11000000000001000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000001000101000111101011100", b"00111110111100001010001111011000"), -- -2.07 + 2.54 = 0.47
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100011110101110000101", b"10111111100010100011110101110000"), -- 2.7 + -3.78 = -1.08
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111011010111000010100011110"), -- -0.48 + 1.4 = 0.92
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011000010100011110101110", b"00111111100111000010100011110101"), -- 2.1 + -0.88 = 1.22
	(b"01000000001010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111110101111010111000010100100", b"01000000000100010100011110101110"), -- 2.64 + -0.37 = 2.27
	(b"11000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000001000111101011100001010", b"00111101010011001100110011000000"), -- -2.51 + 2.56 = 0.05
	(b"00111111111001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000001011000010100011110110", b"01000000100100000000000000000000"), -- 1.81 + 2.69 = 4.5
	(b"11000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111110001111010111000010100", b"10111111010111000010100011111000"), -- -2.42 + 1.56 = -0.86
	(b"11000000000011101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111111001111010111000010100", b"11000000100000010100011110101110"), -- -2.23 + -1.81 = -4.04
	(b"01000000000110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111110100011110101110000110000"), -- 2.38 + -2.1 = 0.28
	(b"01000000000101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111110100001010001111010111", b"00111111001110101110000101000110"), -- 2.36 + -1.63 = 0.73
	(b"01000000000101111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"01000000010100000000000000000000"), -- 2.37 + 0.88 = 3.25
	(b"00111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111100100011110101110000101", b"10111111010001111010111000010100"), -- 0.36 + -1.14 = -0.78
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111110010011001100110011010000"), -- -2.7 + 2.5 = -0.2
	(b"01000000000101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110001111010111000010100", b"01000000011110100011110101110000"), -- 2.35 + 1.56 = 3.91
	(b"01000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110011101011100001010001111", b"01000000010000111101011100001010"), -- 2.82 + 0.24 = 3.06
	(b"11000000000101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111111111101011100001010010", b"11000000100010011110101110000101"), -- -2.32 + -1.99 = -4.31
	(b"00111111100110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111100111010111000010100100", b"01000000000111000010100011110110"), -- 1.21 + 1.23 = 2.44
	(b"01000000000001000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000000010111000010100011111", b"10111101111000010100011111000000"), -- 2.07 + -2.18 = -0.11
	(b"00111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111110100001010001111010111", b"01000000000010001111010111000010"), -- 0.51 + 1.63 = 2.14
	(b"01000000010011101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000100110101000111101011100"), -- 3.23 + 1.6 = 4.83
	(b"11000000000000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111011101011100001010001111", b"10111111100010100011110101110000"), -- -2.04 + 0.96 = -1.08
	(b"00111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000001011000010100011110110", b"11000000000011001100110011001101"), -- 0.49 + -2.69 = -2.2
	(b"01000000010010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000110100011110101110001", b"01000000101100010100011110101110"), -- 3.13 + 2.41 = 5.54
	(b"10111110110101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000011001010001111010111000", b"11000000100000000000000000000000"), -- -0.42 + -3.58 = -4
	(b"11000000001100011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000000101111010111000010100", b"10111110110100011110101110001000"), -- -2.78 + 2.37 = -0.41
	(b"11000000010000011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000010100000000000000000000", b"00111110011000010100011110110000"), -- -3.03 + 3.25 = 0.22
	(b"11000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111101010111000010100011111", b"11000000100001001100110011001101"), -- -2.81 + -1.34 = -4.15
	(b"01000000000101111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111001000010100011110101110", b"01000000010000000000000000000000"), -- 2.37 + 0.63 = 3
	(b"00111101011101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000011110100011110101110001", b"01000000011111100001010001111011"), -- 0.06 + 3.91 = 3.97
	(b"11000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011001000111101011100001", b"11000000111001001100110011001100"), -- -3.58 + -3.57 = -7.15
	(b"01000000001011100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110101110000101000111101100", b"01000000010001010001111010111000"), -- 2.72 + 0.36 = 3.08
	(b"01000000000101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000010111100001010001111011", b"10111111100011100001010001111100"), -- 2.36 + -3.47 = -1.11
	(b"11000000001001000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000010111100001010001111011", b"11000000110000010100011110101110"), -- -2.57 + -3.47 = -6.04
	(b"10111111111010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000011011010111000010100100", b"00111111111100001010001111010111"), -- -1.83 + 3.71 = 1.88
	(b"10111111110010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000010110101110000101001000", b"00111111111010100011110101110001"), -- -1.59 + 3.42 = 1.83
	(b"01000000011111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000011101110000101000111101", b"01000000111110110011001100110011"), -- 3.99 + 3.86 = 7.85
	(b"00111111111011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000100101010001111010111000"), -- 1.86 + 2.8 = 4.66
	(b"00111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000010101111010111000010100", b"01000000011101100110011001100110"), -- 0.48 + 3.37 = 3.85
	(b"11000000010111110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000000001011100001010001111", b"11000000101100101000111101011100"), -- -3.49 + -2.09 = -5.58
	(b"11000000011010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"10111110111000010100011110110000"), -- -3.64 + 3.2 = -0.44
	(b"10111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000001101010001111010111000", b"11000000010011100001010001111010"), -- -0.39 + -2.83 = -3.22
	(b"01000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000010111100001010001111011", b"10111111100001100110011001100110"), -- 2.42 + -3.47 = -1.05
	(b"10111111110101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000000010000101000111101100", b"11000000011100101000111101011100"), -- -1.66 + -2.13 = -3.79
	(b"10111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000011111010111000010100100", b"01000000011000010100011110101110"), -- -0.44 + 3.96 = 3.52
	(b"10111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111101001010001111010111000"), -- -0.34 + -0.95 = -1.29
	(b"01000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"01000000011101100110011001100110"), -- 3.01 + 0.84 = 3.85
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111101111101011100001010010", b"11000000000110100011110101110001"), -- -0.92 + -1.49 = -2.41
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000010111010111000010100100", b"01000000001001100110011001100110"), -- -0.86 + 3.46 = 2.6
	(b"11000000010011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010101110000101000111101", b"11000000000110011001100110011010"), -- -3.24 + 0.84 = -2.4
	(b"11000000010110100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010101110000101000111101", b"10111101010011001100110100000000"), -- -3.41 + 3.36 = -0.0500002
	(b"00111111101111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000010011000010100011110110", b"10111111110111000010100011110110"), -- 1.47 + -3.19 = -1.72
	(b"11000000001101010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000000010100011110101110001", b"10111111001010111000010100011100"), -- -2.83 + 2.16 = -0.67
	(b"01000000001001000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111110111010111000010100100", b"01000000100010011001100110011010"), -- 2.57 + 1.73 = 4.3
	(b"01000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000001011100001010001111011"), -- 2.42 + 0.3 = 2.72
	(b"10111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110111110101110000101001000", b"00111110110100011110101110000110"), -- -0.08 + 0.49 = 0.41
	(b"10111111110111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000100011011100001010010000"), -- -1.73 + -2.7 = -4.43
	(b"11000000011001110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111000111101011100001010010", b"11000000100001110101110000101001"), -- -3.61 + -0.62 = -4.23
	(b"11000000001110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"11000000011110000101000111101100"), -- -2.92 + -0.96 = -3.88
	(b"11000000010010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000000100111101011100001010", b"11000000101011110000101000111110"), -- -3.16 + -2.31 = -5.47
	(b"01000000000010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000010110000101000111101100", b"10111111100111000010100011110110"), -- 2.16 + -3.38 = -1.22
	(b"01000000000101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000000000010100011110101110"), -- 2.32 + -0.3 = 2.02
	(b"10111111111010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111101111101011100001010010", b"11000000010101010001111010111000"), -- -1.84 + -1.49 = -3.33
	(b"00111111101110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000001111101011100001010010", b"10111111110001010001111010111000"), -- 1.44 + -2.98 = -1.54
	(b"11000000000001110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111110100110011001100110011", b"10111110111010111000010100011100"), -- -2.11 + 1.65 = -0.46
	(b"01000000000001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000001100000000000000000000", b"01000000100110101000111101011100"), -- 2.08 + 2.75 = 4.83
	(b"00111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111000001111010111000010100", b"00111111011111010111000010100100"), -- 0.46 + 0.53 = 0.99
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"01000000011011000010100011110110"), -- 3.7 + -0.01 = 3.69
	(b"10111111101110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111101010100011110101110001", b"11000000001100010100011110101110"), -- -1.44 + -1.33 = -2.77
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000001100011110101110000101", b"00111111111011100001010001111010"), -- -0.92 + 2.78 = 1.86
	(b"00111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111011000111101011100001010"), -- 0.99 + -0.1 = 0.89
	(b"11000000010110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000010001111010111000010100", b"11000000110100011001100110011010"), -- -3.43 + -3.12 = -6.55
	(b"01000000010001000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110001000111101011100001010", b"01000000010011101011100001010010"), -- 3.07 + 0.16 = 3.23
	(b"11000000000110111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010001111010111000010100", b"10111111110100110011001100110100"), -- -2.43 + 0.78 = -1.65
	(b"01000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111010000101000111101011100", b"01000000000000110011001100110011"), -- 2.81 + -0.76 = 2.05
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111110100011110101110000101001", b"00111110000110011001100110011010"), -- 0.43 + -0.28 = 0.15
	(b"11000000011100101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111111001111010111000010100", b"10111111111111010111000010100100"), -- -3.79 + 1.81 = -1.98
	(b"01000000011010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011110101110000101001", b"10111101101110000101000111100000"), -- 3.65 + -3.74 = -0.0899999
	(b"00111111111111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111110011110101110000101001", b"00111110101111010111000010100100"), -- 1.99 + -1.62 = 0.37
	(b"01000000000000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111111001010001111010111000", b"00111110011000010100011110110000"), -- 2.01 + -1.79 = 0.22
	(b"01000000011010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110101011100001010001111", b"01000000101010100011110101110001"), -- 3.65 + 1.67 = 5.32
	(b"00111110111000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000000101110000101000111101", b"01000000001100110011001100110011"), -- 0.44 + 2.36 = 2.8
	(b"10111111111000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000000010101110000101001000", b"11000000011111000010100011110110"), -- -1.77 + -2.17 = -3.94
	(b"00111111100101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000011110111000010100011111", b"01000000101000101110000101001000"), -- 1.16 + 3.93 = 5.09
	(b"11000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111110010001111010111000011", b"11000000100011000111101011100001"), -- -2.82 + -1.57 = -4.39
	(b"01000000000001000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000010011010111000010100100", b"01000000101010001111010111000010"), -- 2.07 + 3.21 = 5.28
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000100001001100110011001101"), -- -0.65 + -3.5 = -4.15
	(b"11000000010011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000000000110011001100110011", b"10111111100101011100001010010000"), -- -3.22 + 2.05 = -1.17
	(b"10111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000000000001010001111010111", b"00111111100110011001100110011010"), -- -0.81 + 2.01 = 1.2
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111100001000111101011100001010", b"10111101010011001100110011001100"), -- -0.04 + -0.01 = -0.05
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000000011010111000010100100"), -- -0.79 + 3 = 2.21
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110000101000111101100", b"01000000111100101000111101011100"), -- 3.7 + 3.88 = 7.58
	(b"01000000001101010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111100010001111010111000100"), -- 2.83 + -3.9 = -1.07
	(b"01000000010001000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000101110111101011100001010"), -- 3.07 + 2.8 = 5.87
	(b"00111111111000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"00111111111101000111101011100001"), -- 1.78 + 0.13 = 1.91
	(b"11000000011101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111110100110011001100110011", b"11000000101100000101000111101011"), -- -3.86 + -1.65 = -5.51
	(b"11000000011100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111111101110000101000111101", b"11000000101101111010111000010100"), -- -3.81 + -1.93 = -5.74
	(b"01000000011101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001000111101011100001010", b"01000000010011010111000010100100"), -- 3.85 + -0.64 = 3.21
	(b"11000000001011010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000000111100001010001111011", b"11000000101001011100001010010000"), -- -2.71 + -2.47 = -5.18
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011010100011110101110001", b"11000000110010111000010100011111"), -- -2.7 + -3.66 = -6.36
	(b"01000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101111011100001010010000"), -- 2.93 + 3 = 5.93
	(b"01000000010001011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111100110000101000111101100", b"01000000100010001111010111000010"), -- 3.09 + 1.19 = 4.28
	(b"00111111110100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111100111010111000010100100", b"00111110110100011110101110000100"), -- 1.64 + -1.23 = 0.41
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111111010111000010100100", b"00111111011110101110000101001000"), -- -1 + 1.98 = 0.98
	(b"01000000010010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000010000011110101110000101", b"01000000110001010001111010111000"), -- 3.13 + 3.03 = 6.16
	(b"00111111111011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111101101000111101011100001010", b"00111111111000111101011100001010"), -- 1.86 + -0.08 = 1.78
	(b"11000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000001001000111101011100001", b"11000000110100011001100110011010"), -- -3.98 + -2.57 = -6.55
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000001110100011110101110000"), -- 0.81 + 2.1 = 2.91
	(b"00111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111111011001100110011001101", b"01000000001100010100011110101110"), -- 0.92 + 1.85 = 2.77
	(b"10111110101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"10111101010011001100110011010000"), -- -0.36 + 0.31 = -0.05
	(b"11000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000000111101011100001010010", b"11000000100111110000101000111110"), -- -2.49 + -2.48 = -4.97
	(b"01000000010111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000010101100110011001100110", b"01000000110110010100011110101110"), -- 3.44 + 3.35 = 6.79
	(b"01000000001101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000000000010100011110101110", b"01000000100110111000010100011110"), -- 2.84 + 2.02 = 4.86
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110101011100001010001111", b"10111110101111010111000010100100"), -- 1.3 + -1.67 = -0.37
	(b"00111111100011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111101111000010100011110110", b"10111110101110000101000111101100"), -- 1.11 + -1.47 = -0.36
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110000110011001100110011010", b"11000000000100000000000000000000"), -- -2.1 + -0.15 = -2.25
	(b"00111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011111000010100011110110"), -- 0.64 + 3.3 = 3.94
	(b"00111111111000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000001000010100011110101110", b"01000000100010001111010111000010"), -- 1.76 + 2.52 = 4.28
	(b"11000000011010000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111100111000010100011110110", b"11000000100110110011001100110100"), -- -3.63 + -1.22 = -4.85
	(b"00111111111111000010100011110110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111111011110101110000101001"), -- 1.97 + -0.1 = 1.87
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000000100101000111101011100", b"00111111111101011100001010001111"), -- -0.37 + 2.29 = 1.92
	(b"01000000000010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000011111001100110011001101", b"10111111111001010001111010111000"), -- 2.16 + -3.95 = -1.79
	(b"10111111100000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000011100000000000000000000", b"01000000001011100001010001111011"), -- -1.03 + 3.75 = 2.72
	(b"00111111110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111110100110011001100110011", b"01000000010101111010111000010100"), -- 1.72 + 1.65 = 3.37
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011010001111010111000011", b"00111110100001010001111010111010"), -- -0.65 + 0.91 = 0.26
	(b"01000000001011000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000011111010111000010100100", b"01000000110101001100110011001101"), -- 2.69 + 3.96 = 6.65
	(b"10111111011100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111101000010100011110101110"), -- -0.94 + 2.2 = 1.26
	(b"01000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000000011110101110000101001", b"00111111101010111000010100011110"), -- 3.58 + -2.24 = 1.34
	(b"10111111110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111110101011100001010001111", b"00111100111101011100001010000000"), -- -1.64 + 1.67 = 0.03
	(b"11000000011111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111101111101011100001010010", b"11000000000111100001010001111011"), -- -3.96 + 1.49 = -2.47
	(b"10111111100101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111000011001100110011001101", b"10111111000111101011100001010001"), -- -1.17 + 0.55 = -0.62
	(b"01000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000001010101110000101001000", b"00111110000110011001100110010000"), -- 2.82 + -2.67 = 0.15
	(b"01000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111001011100001010001111011", b"01000000010010101110000101001000"), -- 2.49 + 0.68 = 3.17
	(b"00111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000111101011100001010", b"00111111100010100011110101110000"), -- 0.05 + 1.03 = 1.08
	(b"11000000000111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"11000000010110011001100110011010"), -- -2.45 + -0.95 = -3.4
	(b"10111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000011011101011100001010010", b"11000000100100111101011100001010"), -- -0.89 + -3.73 = -4.62
	(b"00111111111001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"00111111101011001100110011001100"), -- 1.79 + -0.44 = 1.35
	(b"10111111101101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111100101000111101011100001", b"10111110100010100011110101110000"), -- -1.43 + 1.16 = -0.27
	(b"11000000011000011110101110000101", b"00000000000000000000000000000000"),
	(b"00111110001110000101000111101100", b"11000000010101100110011001100110"), -- -3.53 + 0.18 = -3.35
	(b"11000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"00111110101100110011001100110011", b"11000000001001010001111010111001"), -- -2.93 + 0.35 = -2.58
	(b"11000000000110100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"10111111110011110101110000101010"), -- -2.41 + 0.79 = -1.62
	(b"10111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010110101110000101001000", b"01000000001010000101000111101100"), -- -0.79 + 3.42 = 2.63
	(b"10111111111101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111111111010111000010100100", b"00111101100011110101110000110000"), -- -1.91 + 1.98 = 0.0700001
	(b"11000000011111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011010100011110101110001", b"11000000111100111000010100011111"), -- -3.95 + -3.66 = -7.61
	(b"01000000001111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000010100011110101110", b"00111110110111000010100011111000"), -- 2.95 + -2.52 = 0.43
	(b"00111111101111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000000001011100001010001111", b"10111111000111000010100011110100"), -- 1.48 + -2.09 = -0.61
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000011101111010111000010100", b"01000000010001011100001010001111"), -- -0.78 + 3.87 = 3.09
	(b"11000000000110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111111111101011100001010010", b"11000000100010111101011100001010"), -- -2.38 + -1.99 = -4.37
	(b"01000000010101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001011100001010001111", b"10111110011101011100001010010000"), -- 3.35 + -3.59 = -0.24
	(b"10111111111101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111101101000111101011100001", b"11000000010101000111101011100001"), -- -1.91 + -1.41 = -3.32
	(b"01000000011000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000001000011110101110000101", b"01000000110000011001100110011010"), -- 3.52 + 2.53 = 6.05
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011110101110000101001000", b"01000000001100011110101110000101"), -- 1.8 + 0.98 = 2.78
	(b"10111110111110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111110000010100011110101110", b"11000000000000000000000000000000"), -- -0.49 + -1.51 = -2
	(b"11000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000011101011100001010001111", b"00111111100000111101011100001010"), -- -2.81 + 3.84 = 1.03
	(b"00111111101111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000000110000101000111101100", b"01000000011101110000101000111110"), -- 1.48 + 2.38 = 3.86
	(b"00111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111110000101000111101011100", b"01000000000010011001100110011010"), -- 0.63 + 1.52 = 2.15
	(b"01000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111101100001010001111010111", b"00111111101101110000101000111101"), -- 2.81 + -1.38 = 1.43
	(b"11000000001010101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111100000101000111101011100", b"11000000011011000010100011110110"), -- -2.67 + -1.02 = -3.69
	(b"00111111110110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111100110101110000101001000", b"01000000001110011001100110011010"), -- 1.69 + 1.21 = 2.9
	(b"01000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111111000001010001111010111000", b"01000000010000011110101110000101"), -- 2.51 + 0.52 = 3.03
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111110110011001100110011001100"), -- 1.6 + -2 = -0.4
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111111010111000010100100", b"10111101111101011100001010000000"), -- -2.1 + 1.98 = -0.12
	(b"10111111010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110111100001010001111010111", b"10111110100011110101110000101001"), -- -0.75 + 0.47 = -0.28
	(b"01000000000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010011000010100011110110", b"01000000101001111010111000010100"), -- 2.05 + 3.19 = 5.24
	(b"00111101101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"00111111011101011100001010001111"), -- 0.08 + 0.88 = 0.96
	(b"11000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111110001111010111000010100", b"11000000100000100011110101110000"), -- -2.51 + -1.56 = -4.07
	(b"11000000010100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000010111001100110011001101", b"00111110010000101000111101100000"), -- -3.26 + 3.45 = 0.19
	(b"10111111101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111110010100011110101110001", b"00111110000011110101110000101000"), -- -1.44 + 1.58 = 0.14
	(b"10111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111111101110000101000111101", b"11000000010111110101110000101000"), -- -1.56 + -1.93 = -3.49
	(b"01000000000011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000011110101110000101001000", b"10111111110110011001100110011010"), -- 2.22 + -3.92 = -1.7
	(b"10111111101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111101110011001100110011010", b"00111100001000111101011100000000"), -- -1.44 + 1.45 = 0.00999999
	(b"10111111110110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111111011001100110011001101", b"11000000011000111101011100001010"), -- -1.71 + -1.85 = -3.56
	(b"00111111100010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"00111110100000000000000000000010"), -- 1.07 + -0.82 = 0.25
	(b"01000000011001110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000010010000101000111101100", b"00111110111101011100001010001000"), -- 3.61 + -3.13 = 0.48
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111101000000000000000000000", b"00111111110010001111010111000010"), -- 0.32 + 1.25 = 1.57
	(b"00111110110111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000001110111000010100011111", b"01000000010101110000101000111110"), -- 0.43 + 2.93 = 3.36
	(b"10111111100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001010111000010100011111", b"11000000011101010001111010111000"), -- -1.15 + -2.68 = -3.83
	(b"10111111100001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000000000001010001111010111", b"11000000010000110011001100110011"), -- -1.04 + -2.01 = -3.05
	(b"01000000001111110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000010001000111101011100001", b"10111101101000111101011100000000"), -- 2.99 + -3.07 = -0.0799999
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001000111101011100001", b"10111101100011110101110000100000"), -- 3.5 + -3.57 = -0.0699999
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111101100011110101110000101", b"10111111100010001111010111000010"), -- 0.32 + -1.39 = -1.07
	(b"00111111110100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111110111010111000010100011111", b"00111111100101011100001010001111"), -- 1.63 + -0.46 = 1.17
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111101001010001111010111000", b"00111111110101011100001010001111"), -- 0.38 + 1.29 = 1.67
	(b"11000000010001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111100001111010111000010100", b"11000000100001011100001010001111"), -- -3.12 + -1.06 = -4.18
	(b"11000000000100101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000000111110101110000101001", b"00111110010011001100110011010000"), -- -2.29 + 2.49 = 0.2
	(b"10111111000001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111010100011110101110000101", b"00111110100101000111101011100010"), -- -0.53 + 0.82 = 0.29
	(b"00111111000010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000011111100001010001111011", b"11000000010110111000010100011111"), -- 0.54 + -3.97 = -3.43
	(b"00111111000001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111111101110000101000111101", b"10111111101101000111101011100001"), -- 0.52 + -1.93 = -1.41
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011000010100011110110", b"10111111111111101011100001010010"), -- 1.2 + -3.19 = -1.99
	(b"00111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111010000000000000000000000"), -- 0.55 + 0.2 = 0.75
	(b"00111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000001011110101110000101001", b"01000000001111100001010001111011"), -- 0.23 + 2.74 = 2.97
	(b"00111111111100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111111000000000000000000000", b"00111110000011110101110000101000"), -- 1.89 + -1.75 = 0.14
	(b"01000000001001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000000010000101000111101100", b"01000000100110000000000000000000"), -- 2.62 + 2.13 = 4.75
	(b"01000000001010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"01000000001110111000010100011111"), -- 2.68 + 0.25 = 2.93
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000010010100011110101110001", b"11000000011111101011100001010010"), -- -0.82 + -3.16 = -3.98
	(b"10111111101011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110101110000101001000", b"11000000010000111101011100001010"), -- -1.35 + -1.71 = -3.06
	(b"10111111100111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111110001000111101011100001010", b"10111111101100011110101110000101"), -- -1.23 + -0.16 = -1.39
	(b"10111111011110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000111010111000010100100", b"00111111101111101011100001010010"), -- -0.97 + 2.46 = 1.49
	(b"11000000000101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110100011110101110000101", b"11000000001100001010001111010111"), -- -2.35 + -0.41 = -2.76
	(b"00111111111000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110111010111000010100100", b"01000000010111101011100001010010"), -- 1.75 + 1.73 = 3.48
	(b"01000000011000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000010111010111000010100100", b"00111101110011001100110011000000"), -- 3.56 + -3.46 = 0.0999999
	(b"01000000000010101110000101001000", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"01000000000011010111000010100100"), -- 2.17 + 0.04 = 2.21
	(b"01000000000101010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000010100000000000000000000", b"01000000101100101000111101011100"), -- 2.33 + 3.25 = 5.58
	(b"01000000001101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111111010111000010100011110100"), -- 2.86 + -2 = 0.86
	(b"11000000011101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"10111110100001010001111010111000"), -- -3.86 + 3.6 = -0.26
	(b"00111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111101000010100011110101110", b"01000000001101000111101011100001"), -- 1.56 + 1.26 = 2.82
	(b"00111111111010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000011110000101000111101100", b"01000000101101100110011001100111"), -- 1.82 + 3.88 = 5.7
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000101000111101011100", b"10111110011000010100011110101100"), -- 0.8 + -1.02 = -0.22
	(b"10111111001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"10111111010011110101110000101001"), -- -0.64 + -0.17 = -0.81
	(b"00111111011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100001010001111010111", b"11000000000100111101011100001010"), -- 0.95 + -3.26 = -2.31
	(b"01000000001000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000010110001111010111000011", b"10111111010101000111101011100100"), -- 2.56 + -3.39 = -0.83
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001100001010001111010111", b"01000000001100010100011110101110"), -- 0.01 + 2.76 = 2.77
	(b"11000000010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000000100011110101110000101"), -- -3.28 + 1 = -2.28
	(b"10111111110011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000010101000111101011100010"), -- -1.62 + -1.7 = -3.32
	(b"11000000011101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111110010111000010100011111", b"11000000000100010100011110101110"), -- -3.86 + 1.59 = -2.27
	(b"01000000000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000101000111101011100", b"01000000100101100001010001111011"), -- 2.15 + 2.54 = 4.69
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000001100000000000000000000", b"11000000010111000010100011110110"), -- -0.69 + -2.75 = -3.44
	(b"01000000010111110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110111110101110000101001000", b"01000000010000000000000000000000"), -- 3.49 + -0.49 = 3
	(b"11000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000011100111101011100001010", b"11000000110010100011110101110000"), -- -2.51 + -3.81 = -6.32
	(b"11000000011000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"10111111011100110011001100110100"), -- -3.55 + 2.6 = -0.95
	(b"10111111101100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000011000011110101110000101", b"11000000100111010111000010100100"), -- -1.39 + -3.53 = -4.92
	(b"11000000001110100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111100010100011110101110001", b"11000000011111110101110000101010"), -- -2.91 + -1.08 = -3.99
	(b"01000000011010101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000001000110011001100110011", b"01000000110001110000101000111110"), -- 3.67 + 2.55 = 6.22
	(b"11000000010101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011111001100110011001101", b"11000000111010011001100110011010"), -- -3.35 + -3.95 = -7.3
	(b"01000000010010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110100001010001111010111", b"01000000100110001111010111000011"), -- 3.15 + 1.63 = 4.78
	(b"01000000000010101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"01000000001101000111101011100010"), -- 2.17 + 0.65 = 2.82
	(b"01000000001100101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111111101011100001010001111", b"01000000100101101011100001010010"), -- 2.79 + 1.92 = 4.71
	(b"10111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111100011100001010001111011", b"00111110100101000111101011100010"), -- -0.82 + 1.11 = 0.29
	(b"11000000011000011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111110110000101000111101100", b"10111111111010111000010100011110"), -- -3.53 + 1.69 = -1.84
	(b"11000000010001011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000001011000010100011110110", b"11000000101110001111010111000010"), -- -3.09 + -2.69 = -5.78
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001101110000101000111101", b"01000000011100000000000000000000"), -- 0.89 + 2.86 = 3.75
	(b"01000000010100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000001010000101000111101100", b"00111111001001100110011001100100"), -- 3.28 + -2.63 = 0.65
	(b"11000000001001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010000011110101110000101", b"11000000101101001100110011001100"), -- -2.62 + -3.03 = -5.65
	(b"10111111110110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111101100011110101110000101", b"10111110101000111101011100001100"), -- -1.71 + 1.39 = -0.32
	(b"01000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"01000000010100101000111101011100"), -- 3.01 + 0.28 = 3.29
	(b"01000000010110111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000001101011100001010001111", b"01000000110010001010001111010111"), -- 3.43 + 2.84 = 6.27
	(b"01000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111101000111101011100001010", b"01000000000100110011001100110011"), -- 3.58 + -1.28 = 2.3
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"10111110110111000010100011110111"), -- -0.72 + 0.29 = -0.43
	(b"00111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000010011000010100011110110", b"11000000010000011110101110000101"), -- 0.16 + -3.19 = -3.03
	(b"00111111100000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000011110000101000111101100", b"11000000001101111010111000010101"), -- 1.01 + -3.88 = -2.87
	(b"00111110001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111101101110000101000111101", b"00111111110011100001010001111010"), -- 0.18 + 1.43 = 1.61
	(b"01000000001110001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000001001111010111000010100", b"01000000101100000101000111101100"), -- 2.89 + 2.62 = 5.51
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000011101011100001010010", b"11000000101000001111010111000010"), -- -2.8 + -2.23 = -5.03
	(b"00111111100101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000100010111101011100001010"), -- 1.17 + 3.2 = 4.37
	(b"11000000001000011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000011100000000000000000000", b"00111111100111000010100011110110"), -- -2.53 + 3.75 = 1.22
	(b"10111111100001100110011001100110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"10111111100001100110011001100110"), -- -1.05 + 0 = -1.05
	(b"10111111100110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111010111000010100011110110", b"10111110101100110011001100110100"), -- -1.21 + 0.86 = -0.35
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010011000010100011110110", b"01000000010111010111000010100100"), -- 0.27 + 3.19 = 3.46
	(b"01000000001111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111100101110000101000111101", b"01000000100001010001111010111000"), -- 2.98 + 1.18 = 4.16
	(b"00111111111100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"00111111101001100110011001100110"), -- 1.89 + -0.59 = 1.3
	(b"11000000011000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000001000001010001111010111", b"11000000110000011001100110011010"), -- -3.54 + -2.51 = -6.05
	(b"11000000000100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111110111101011100001010010", b"10111111000010100011110101110000"), -- -2.28 + 1.74 = -0.54
	(b"11000000000100101000111101011100", b"00000000000000000000000000000000"),
	(b"00111110100011110101110000101001", b"11000000000000001010001111010111"), -- -2.29 + 0.28 = -2.01
	(b"11000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000011101000111101011100001", b"10111101011101011100001011000000"), -- -3.88 + 3.82 = -0.0600002
	(b"01000000000010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000000011110101110000101", b"01000000100001010001111010111000"), -- 2.13 + 2.03 = 4.16
	(b"11000000001011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000010111000010100011110110", b"00111111001110000101000111101100"), -- -2.72 + 3.44 = 0.72
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110111101011100001010010", b"11000000101100010100011110101110"), -- -3.8 + -1.74 = -5.54
	(b"11000000011110111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111111101011100001010001111", b"11000000101110110011001100110011"), -- -3.93 + -1.92 = -5.85
	(b"00111111101010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000000111101011100001010010"), -- 1.32 + -3.8 = -2.48
	(b"11000000011001000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000000000101000111101011100", b"10111111110000111101011100001010"), -- -3.57 + 2.04 = -1.53
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110011010111000010100011111", b"10111111000100011110101110000101"), -- -0.8 + 0.23 = -0.57
	(b"10111111110101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000101010001111010111000010"), -- -1.68 + -3.6 = -5.28
	(b"10111111111000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111111110011001100110011010", b"00111110010000101000111101100000"), -- -1.76 + 1.95 = 0.19
	(b"00111111111010111000010100011111", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"01000000000001011100001010010000"), -- 1.84 + 0.25 = 2.09
	(b"01000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000000001011100001010001111", b"01000000101000001010001111010111"), -- 2.93 + 2.09 = 5.02
	(b"01000000010100010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"00111111110010001111010111000010"), -- 3.27 + -1.7 = 1.57
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110001111010111000011", b"11000000010110001111010111000011"), -- -1 + -2.39 = -3.39
	(b"00111110110001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000001011000010100011110110", b"01000000010001010001111010111000"), -- 0.39 + 2.69 = 3.08
	(b"11000000000111100001010001111011", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"11000000001000000000000000000000"), -- -2.47 + -0.03 = -2.5
	(b"10111111001100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000000001010001111010111000", b"11000000001100010100011110101110"), -- -0.69 + -2.08 = -2.77
	(b"00111111110010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000100001100001010001111011"), -- 1.59 + 2.6 = 4.19
	(b"11000000000010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000000111001100110011001101", b"11000000100101000010100011110110"), -- -2.18 + -2.45 = -4.63
	(b"10111101001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111101000000000000000000000", b"10111111101001010001111010111000"), -- -0.04 + -1.25 = -1.29
	(b"10111111010001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000001010101110000101001000"), -- -0.77 + -1.9 = -2.67
	(b"01000000011000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000011000010100011110101110", b"01000000111000011110101110000101"), -- 3.54 + 3.52 = 7.06
	(b"11000000001110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000011110000101000111101100", b"00111111011101011100001010010000"), -- -2.92 + 3.88 = 0.96
	(b"11000000011111100001010001111011", b"00000000000000000000000000000000"),
	(b"00111111110001100110011001100110", b"11000000000110101110000101001000"), -- -3.97 + 1.55 = -2.42
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000110000101000111101100", b"00111111100010100011110101110010"), -- -1.3 + 2.38 = 1.08
	(b"00111111100010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000010011100001010001111011", b"01000000100010010100011110101110"), -- 1.07 + 3.22 = 4.29
	(b"01000000010111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011101011100001010010", b"01000000111001011100001010010000"), -- 3.45 + 3.73 = 7.18
	(b"11000000001011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000000110101110000101001000", b"11000000101001010001111010111000"), -- -2.74 + -2.42 = -5.16
	(b"10111111000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001111010111000010100", b"11000000000101110000101000111101"), -- -0.55 + -1.81 = -2.36
	(b"10111111100111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111110100111101011100001010010", b"10111111011011100001010001111011"), -- -1.24 + 0.31 = -0.93
	(b"10111111101110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111010110011001100110011010"), -- -1.45 + 0.6 = -0.85
	(b"11000000011101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000111011010111000010100100"), -- -3.82 + -3.6 = -7.42
	(b"10111111111011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000011101110000101000111101", b"11000000101101110101110000101001"), -- -1.87 + -3.86 = -5.73
	(b"01000000010001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000000101000111101011100001", b"01000000101011100001010001111010"), -- 3.12 + 2.32 = 5.44
	(b"00111111110010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111101101000111101011100001", b"00111110001110000101000111110000"), -- 1.59 + -1.41 = 0.18
	(b"11000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000110001010111000010100100"), -- -2.97 + -3.2 = -6.17
	(b"00111111111110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111010100011110101110000101", b"01000000001100001010001111010111"), -- 1.94 + 0.82 = 2.76
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100001010001111010111000", b"00111111101001010001111010111000"), -- 0.25 + 1.04 = 1.29
	(b"10111110011101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000011001010001111010111000", b"01000000010101011100001010001111"), -- -0.24 + 3.58 = 3.34
	(b"10111111011111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"10111111101101110000101000111110"), -- -0.99 + -0.44 = -1.43
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110101100110011001100110011", b"01000000001010011001100110011001"), -- 2.3 + 0.35 = 2.65
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010001111010111000010100", b"00111111111100001010001111010111"), -- 1.1 + 0.78 = 1.88
	(b"10111111111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111111100001010001111010111", b"10111101001000111101011100000000"), -- -1.92 + 1.88 = -0.04
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011110101110000101001", b"11000000000000010100011110101110"), -- -0.4 + -1.62 = -2.02
	(b"01000000011111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000101111010111000010100", b"00111111110010100011110101110010"), -- 3.95 + -2.37 = 1.58
	(b"01000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000001011101011100001010010", b"01000000101001001100110011001101"), -- 2.42 + 2.73 = 5.15
	(b"10111111011101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111110101000111101011100001"), -- -0.96 + -0.7 = -1.66
	(b"11000000000101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000001001110000101000111101", b"00111110100000000000000000000000"), -- -2.36 + 2.61 = 0.25
	(b"10111111111111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111101010001111010111000011", b"11000000010100110011001100110100"), -- -1.98 + -1.32 = -3.3
	(b"01000000000010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001111010111000010100100", b"00111111101101000111101011100010"), -- 2.15 + -0.74 = 1.41
	(b"01000000011011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000011001000111101011100001", b"01000000111010011110101110000101"), -- 3.74 + 3.57 = 7.31
	(b"00111111100101110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111011000010100011110101110", b"01000000000000111101011100001010"), -- 1.18 + 0.88 = 2.06
	(b"11000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111111000010100011110101110", b"11000000000001111010111000010101"), -- -3.88 + 1.76 = -2.12
	(b"11000000010110100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111100110000101000111101100", b"11000000000011100001010001111011"), -- -3.41 + 1.19 = -2.22
	(b"10111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001010100011110101110001", b"01000000000101011100001010010000"), -- -0.32 + 2.66 = 2.34
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"11000000000101011100001010010000"), -- -2.4 + 0.06 = -2.34
	(b"11000000001101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000101000111101011100", b"11000000100010111101011100001010"), -- -2.85 + -1.52 = -4.37
	(b"11000000010110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111100000101000111101011100", b"11000000100011001100110011001101"), -- -3.38 + -1.02 = -4.4
	(b"00111111000000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111111111010111000010100100", b"01000000000111110101110000101001"), -- 0.51 + 1.98 = 2.49
	(b"11000000010111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000011111010111000010100100", b"00111110111110101110000101001000"), -- -3.47 + 3.96 = 0.49
	(b"11000000000111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000001101011100001010001111", b"11000000101010011110101110000101"), -- -2.47 + -2.84 = -5.31
	(b"01000000011001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111111010001111010111000011", b"00111111111001100110011001100101"), -- 3.62 + -1.82 = 1.8
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110000101000111101100", b"11000000110010001111010111000011"), -- -3.9 + -2.38 = -6.28
	(b"10111111010101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000001010111000010100011111", b"11000000011000010100011110101110"), -- -0.84 + -2.68 = -3.52
	(b"01000000011110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000110000101000111101100", b"01000000110010000101000111101100"), -- 3.88 + 2.38 = 6.26
	(b"11000000011110111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000001000101000111101011100", b"11000000110011110000101000111110"), -- -3.93 + -2.54 = -6.47
	(b"01000000011000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"01000000001110111000010100011111"), -- 3.51 + -0.58 = 2.93
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011000111101011100001010", b"00111111010101110000101000111101"), -- -0.05 + 0.89 = 0.84
	(b"11000000011000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111011101011100001010001111", b"11000000100011110101110000101001"), -- -3.52 + -0.96 = -4.48
	(b"01000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000111011110101110000101001"), -- 3.58 + 3.9 = 7.48
	(b"10111111110111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000001000001010001111010111", b"11000000100001111010111000010100"), -- -1.73 + -2.51 = -4.24
	(b"10111111111010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111110000110011001100110011010", b"10111111111111101011100001010010"), -- -1.84 + -0.15 = -1.99
	(b"01000000011011010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111100101110000101000111101", b"01000000100111000111101011100001"), -- 3.71 + 1.18 = 4.89
	(b"10111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010000010100011110101110"), -- -0.38 + 3.4 = 3.02
	(b"01000000010111010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111110011110101110000101001", b"01000000101000101000111101011100"), -- 3.46 + 1.62 = 5.08
	(b"00111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000000111000010100011110110", b"01000000001010100011110101110001"), -- 0.22 + 2.44 = 2.66
	(b"01000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111100001010001111010111000", b"00111111111000101000111101011100"), -- 2.81 + -1.04 = 1.77
	(b"11000000000011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000001101110000101000111101", b"11000000101000110011001100110011"), -- -2.24 + -2.86 = -5.1
	(b"11000000010111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000000000111101011100001010", b"11000000101100000000000000000000"), -- -3.44 + -2.06 = -5.5
	(b"11000000011011101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111111000010100011110101110", b"10111111111111000010100011110110"), -- -3.73 + 1.76 = -1.97
	(b"01000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111110111000010100011110101110", b"01000000001111001100110011001101"), -- 2.51 + 0.44 = 2.95
	(b"11000000000001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000000000110011001100110011", b"11000000100001000010100011110110"), -- -2.08 + -2.05 = -4.13
	(b"11000000001000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000000111110101110000101001", b"10111100111101011100001010000000"), -- -2.52 + 2.49 = -0.03
	(b"11000000001110001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111010101000111101011100001", b"11000000000000111101011100001011"), -- -2.89 + 0.83 = -2.06
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010101100110011001100110", b"10111111001001100110011001100100"), -- 2.7 + -3.35 = -0.65
	(b"11000000011100111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000010111100001010001111011", b"10111110101011100001010001111000"), -- -3.81 + 3.47 = -0.34
	(b"11000000010011000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000010011101011100001010010", b"11000000110011010111000010100100"), -- -3.19 + -3.23 = -6.42
	(b"01000000001101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000000001011100001010001111", b"01000000100111011100001010001111"), -- 2.84 + 2.09 = 4.93
	(b"11000000010011100001010001111011", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"11000000011110100011110101110001"), -- -3.22 + -0.69 = -3.91
	(b"11000000010111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000010101111010111000010100", b"11000000110110110011001100110011"), -- -3.48 + -3.37 = -6.85
	(b"01000000000000011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000011010100011110101110001", b"01000000101101100001010001111011"), -- 2.03 + 3.66 = 5.69
	(b"11000000000101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110110000101000111101100", b"10111111001010001111010111000000"), -- -2.35 + 1.69 = -0.66
	(b"00111111100111000010100011110110", b"00000000000000000000000000000000"),
	(b"11000000011001010001111010111000", b"11000000000101110000101000111101"), -- 1.22 + -3.58 = -2.36
	(b"11000000011111101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000011000110011001100110011", b"10111110110111000010100011111000"), -- -3.98 + 3.55 = -0.43
	(b"11000000010100010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111110111100001010001111011000"), -- -3.27 + 2.8 = -0.47
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011101110000101000111101", b"11000000011010100011110101110000"), -- 0.2 + -3.86 = -3.66
	(b"01000000000000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111000010100011110101110001", b"01000000001001100110011001100110"), -- 2.06 + 0.54 = 2.6
	(b"10111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000000101000111101011100001", b"11000000001001010001111010111000"), -- -0.26 + -2.32 = -2.58
	(b"01000000011010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111110111000010100011110101110", b"01000000010011100001010001111011"), -- 3.66 + -0.44 = 3.22
	(b"10111110011010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000001010000101000111101100", b"11000000001101110000101000111110"), -- -0.23 + -2.63 = -2.86
	(b"10111111110101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000001010000101000111101100", b"00111111011101011100001010010010"), -- -1.67 + 2.63 = 0.96
	(b"00111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"11000000010001111010111000010100", b"11000000000100000000000000000000"), -- 0.87 + -3.12 = -2.25
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000001101100110011001100110", b"11000000001000011110101110000101"), -- 0.32 + -2.85 = -2.53
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111101000111101011100001", b"11000000101100000101000111101011"), -- -3.6 + -1.91 = -5.51
	(b"10111111100010001111010111000011", b"00000000000000000000000000000000"),
	(b"10111110110111000010100011110110", b"10111111110000000000000000000000"), -- -1.07 + -0.43 = -1.5
	(b"10111111110100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111110000111101011100001010", b"10111101111000010100011110110000"), -- -1.64 + 1.53 = -0.11
	(b"00111101111000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111100111101011100001010001111", b"00111101101000111101011100001010"), -- 0.11 + -0.03 = 0.08
	(b"01000000000110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"01000000000000000000000000000000"), -- 2.38 + -0.38 = 2
	(b"10111110100101000111101011100001", b"00000000000000000000000000000000"),
	(b"01000000010001111010111000010100", b"01000000001101010001111010111000"), -- -0.29 + 3.12 = 2.83
	(b"10111111110100001010001111010111", b"00000000000000000000000000000000"),
	(b"01000000001111010111000010100100", b"00111111101010100011110101110001"), -- -1.63 + 2.96 = 1.33
	(b"01000000000001000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111110100001010001111010111", b"01000000011011001100110011001100"), -- 2.07 + 1.63 = 3.7
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111100111101011100001010001111", b"11000000011101111010111000010101"), -- -3.9 + 0.03 = -3.87
	(b"10111111010101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"10111111011000010100011110101110"), -- -0.83 + -0.05 = -0.88
	(b"11000000001100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011000010100011110110", b"10111111000011110101110000101000"), -- -2.75 + 2.19 = -0.56
	(b"01000000010100010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111111011001100110011001101", b"00111111101101011100001010001111"), -- 3.27 + -1.85 = 1.42
	(b"00111110100001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111111101000010100011110101110", b"00111111110000101000111101011100"), -- 0.26 + 1.26 = 1.52
	(b"10111111101000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000011110101110000101001000", b"11000000101001100110011001100110"), -- -1.28 + -3.92 = -5.2
	(b"11000000000010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111100100011110101110000100"), -- -2.16 + 3.3 = 1.14
	(b"01000000001001110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111000001111010111000010100", b"01000000000001010001111010111000"), -- 2.61 + -0.53 = 2.08
	(b"01000000011000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111110000111101011100001010", b"01000000000000001010001111010111"), -- 3.54 + -1.53 = 2.01
	(b"00111111101000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000000000111101011100001010", b"01000000010101010001111010111000"), -- 1.27 + 2.06 = 3.33
	(b"11000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111010011110101110000101001", b"11000000011001111010111000010100"), -- -2.81 + -0.81 = -3.62
	(b"01000000010100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110011101011100001010001111", b"01000000010000001010001111010111"), -- 3.25 + -0.24 = 3.01
	(b"11000000011001110000101000111101", b"00000000000000000000000000000000"),
	(b"00111111101100011110101110000101", b"11000000000011100001010001111010"), -- -3.61 + 1.39 = -2.22
	(b"10111111001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000010101100110011001100110"), -- -0.65 + -2.7 = -3.35
	(b"11000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000010010111000010100011111", b"10111110011101011100001010010000"), -- -3.42 + 3.18 = -0.24
	(b"10111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111010001111010111000010100", b"10111111100011001100110011001100"), -- -0.32 + -0.78 = -1.1
	(b"11000000001111110101110000101001", b"00000000000000000000000000000000"),
	(b"10111110001011100001010001111011", b"11000000010010100011110101110001"), -- -2.99 + -0.17 = -3.16
	(b"10111111111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111111011100110011001100110100"), -- -1.75 + 2.7 = 0.95
	(b"11000000011000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001010001111010111000", b"11000000101010101110000101001000"), -- -3.55 + -1.79 = -5.34
	(b"00111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111000011001100110011001101", b"10111111000010100011110101110001"), -- 0.01 + -0.55 = -0.54
	(b"01000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000001010100011110101110001", b"00111110101100110011001100110000"), -- 3.01 + -2.66 = 0.35
	(b"01000000001100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111111001010001111010111000", b"01000000100100100011110101110000"), -- 2.78 + 1.79 = 4.57
	(b"11000000010011000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000011011000010100011110110"), -- -3.19 + -0.5 = -3.69
	(b"10111111011000010100011110101110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000000001111010111000010100"), -- -0.88 + 3 = 2.12
	(b"11000000001010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111111011100001010001111010100"), -- -2.66 + 3.6 = 0.94
	(b"10111111001000010100011110101110", b"00000000000000000000000000000000"),
	(b"10111111111001111010111000010100", b"11000000000111000010100011110110"), -- -0.63 + -1.81 = -2.44
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110100011110101110000101", b"11000000000011000010100011110101"), -- -2.6 + 0.41 = -2.19
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111001010111000010100011111", b"01000000100011110000101000111101"), -- 3.8 + 0.67 = 4.47
	(b"11000000011110100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000000011000010100011110110", b"10111111110111000010100011110110"), -- -3.91 + 2.19 = -1.72
	(b"01000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111111101000111101011100001", b"00111111100011001100110011001101"), -- 3.01 + -1.91 = 1.1
	(b"11000000000000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111111011011100001010001111011", b"11000000001111110101110000101001"), -- -2.06 + -0.93 = -2.99
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010101010001111010111000", b"01000000101001110101110000101001"), -- 1.9 + 3.33 = 5.23
	(b"11000000011100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"11000000010010000101000111101100"), -- -3.75 + 0.62 = -3.13
	(b"01000000000010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000010101110000101001000", b"01000000100010011001100110011010"), -- 2.13 + 2.17 = 4.3
	(b"11000000001000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"11000000001001011100001010001111"), -- -2.54 + -0.05 = -2.59
	(b"10111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110001110000101000111101100", b"10111111100000111101011100001010"), -- -0.85 + -0.18 = -1.03
	(b"01000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000000110111000010100011111", b"00111101011101011100001010000000"), -- 2.49 + -2.43 = 0.0599999
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000010011100001010001111011", b"11000000000110111000010100011111"), -- 0.79 + -3.22 = -2.43
	(b"01000000011010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111111000111101011100001010", b"00111111111100110011001100110100"), -- 3.68 + -1.78 = 1.9
	(b"11000000000010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000011010111000010100011111", b"00111111110001100110011001100110"), -- -2.13 + 3.68 = 1.55
	(b"01000000000001011100001010001111", b"00000000000000000000000000000000"),
	(b"10111110011010111000010100011111", b"00111111111011100001010001111010"), -- 2.09 + -0.23 = 1.86
	(b"11000000010000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000000000010100011110101110", b"11000000101000001111010111000010"), -- -3.01 + -2.02 = -5.03
	(b"11000000010101111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000001111101011100001010010", b"10111110110001111010111000010000"), -- -3.37 + 2.98 = -0.39
	(b"10111111110111010111000010100100", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"10111111110111010111000010100100"), -- -1.73 + 0 = -1.73
	(b"00111111110011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111011111010111000010100100", b"00111111001000010100011110101110"), -- 1.62 + -0.99 = 0.63
	(b"11000000000001011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111010100011110101110000101", b"11000000001110100011110101110000"), -- -2.09 + -0.82 = -2.91
	(b"10111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000010000001010001111010111", b"01000000000100101000111101011100"), -- -0.72 + 3.01 = 2.29
	(b"11000000010001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"10111101101000111101011100000000"), -- -3.08 + 3 = -0.0799999
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000000010101110000101001000", b"11000000000101010001111010111001"), -- -0.16 + -2.17 = -2.33
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011101111010111000010100", b"01000000111011110000101000111101"), -- 3.6 + 3.87 = 7.47
	(b"11000000001110111000010100011111", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"11000000000010001111010111000011"), -- -2.93 + 0.79 = -2.14
	(b"11000000010111110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111100100011110101110000101", b"11000000100101000010100011110110"), -- -3.49 + -1.14 = -4.63
	(b"01000000000010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000010001000111101011100001", b"01000000101010000000000000000000"), -- 2.18 + 3.07 = 5.25
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010101000111101011100001", b"00111111110111000010100011110101"), -- -1.6 + 3.32 = 1.72
	(b"00111111100101000111101011100001", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000000010001111010111000010"), -- 1.16 + -3.3 = -2.14
	(b"01000000010110001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000000011101011100001010010", b"01000000101100111101011100001010"), -- 3.39 + 2.23 = 5.62
	(b"01000000010011000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111011110000101000111101100", b"01000000100001010001111010111000"), -- 3.19 + 0.97 = 4.16
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011000010100011110110", b"11000000011111110101110000101001"), -- -1.8 + -2.19 = -3.99
	(b"01000000001001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111110100011110101110000101", b"01000000100010000101000111101011"), -- 2.62 + 1.64 = 4.26
	(b"10111111101000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000001101110000101000111101", b"11000000100000111101011100001010"), -- -1.26 + -2.86 = -4.12
	(b"11000000010111100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000000100001010001111010111", b"11000000101101110101110000101001"), -- -3.47 + -2.26 = -5.73
	(b"11000000010110101110000101001000", b"00000000000000000000000000000000"),
	(b"01000000010110100011110101110001", b"10111100001000111101011100000000"), -- -3.42 + 3.41 = -0.00999999
	(b"10111111111110101110000101001000", b"00000000000000000000000000000000"),
	(b"00111111100100110011001100110011", b"10111111010011110101110000101010"), -- -1.96 + 1.15 = -0.81
	(b"10111111110101000111101011100001", b"00000000000000000000000000000000"),
	(b"10111111111001010001111010111000", b"11000000010111001100110011001100"), -- -1.66 + -1.79 = -3.45
	(b"01000000010101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011110101110000101001", b"01000000100111110000101000111101"), -- 3.35 + 1.62 = 4.97
	(b"01000000010000011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111001000010100011110101100"), -- 3.03 + -2.4 = 0.63
	(b"01000000001101010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000001011010111000010100100", b"01000000101100010100011110101110"), -- 2.83 + 2.71 = 5.54
	(b"11000000011101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000111000010100011110110"), -- -3.84 + 1.4 = -2.44
	(b"11000000000010100011110101110001", b"00000000000000000000000000000000"),
	(b"11000000010110111000010100011111", b"11000000101100101110000101001000"), -- -2.16 + -3.43 = -5.59
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000000010001111010111000011", b"01000000000111101011100001010010"), -- 0.34 + 2.14 = 2.48
	(b"01000000001001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000001101110000101000111101", b"10111110011101011100001010010000"), -- 2.62 + -2.86 = -0.24
	(b"11000000011010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"11000000100000001111010111000011"), -- -3.65 + -0.38 = -4.03
	(b"00111111110101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110001011100001010001111011", b"00111111111010111000010100011110"), -- 1.67 + 0.17 = 1.84
	(b"10111110111101011100001010001111", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111110100011110101110000101000"), -- -0.48 + 0.2 = -0.28
	(b"00111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011010111000010100011111", b"00111111100101011100001010010000"), -- 0.25 + 0.92 = 1.17
	(b"10111110100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000101110000101000111101", b"10111111010101110000101000111101"), -- -0.25 + -0.59 = -0.84
	(b"11000000001011010111000010100100", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"11000000001010101110000101001000"), -- -2.71 + 0.04 = -2.67
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000100110011001100110011010"), -- 1.5 + 3.3 = 4.8
	(b"00111110100010100011110101110001", b"00000000000000000000000000000000"),
	(b"01000000011001000111101011100001", b"01000000011101011100001010001111"), -- 0.27 + 3.57 = 3.84
	(b"11000000001110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000001110001111010111000011", b"11000000101110001010001111011000"), -- -2.88 + -2.89 = -5.77
	(b"00111101101110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111110100000000000000000000000", b"00111110101011100001010001111011"), -- 0.09 + 0.25 = 0.34
	(b"01000000001100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000011100011110101110000101", b"10111111100000101000111101011100"), -- 2.76 + -3.78 = -1.02
	(b"11000000010001011100001010001111", b"00000000000000000000000000000000"),
	(b"11000000010111100001010001111011", b"11000000110100011110101110000101"), -- -3.09 + -3.47 = -6.56
	(b"00111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000001011000010100011110110", b"10111111111011110101110000101010"), -- 0.82 + -2.69 = -1.87
	(b"10111111110111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000010111101011100001010010", b"00111111111000010100011110101110"), -- -1.72 + 3.48 = 1.76
	(b"10111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111110100001010001111010111000", b"10111111111010001111010111000010"), -- -1.56 + -0.26 = -1.82
	(b"00111110101011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000011011000010100011110110", b"11000000010101100110011001100111"), -- 0.34 + -3.69 = -3.35
	(b"11000000010100011110101110000101", b"00000000000000000000000000000000"),
	(b"01000000011110101110000101001000", b"00111111001000111101011100001100"), -- -3.28 + 3.92 = 0.64
	(b"11000000000111110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000001110100011110101110001", b"00111110110101110000101001000000"), -- -2.49 + 2.91 = 0.42
	(b"01000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"00111110000001010001111010111000", b"01000000011011010111000010100100"), -- 3.58 + 0.13 = 3.71
	(b"11000000011100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111100100011110101110000101", b"11000000001010001111010111000010"), -- -3.78 + 1.14 = -2.64
	(b"00111111110111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111000111101011100001010010", b"01000000000101011100001010010000"), -- 1.72 + 0.62 = 2.34
	(b"11000000000001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011110111000010100011111", b"11000000110000000101000111101100"), -- -2.08 + -3.93 = -6.01
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011100110011001100110011", b"10111111000011001100110011001100"), -- 0.4 + -0.95 = -0.55
	(b"10111111100001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000001001000111101011100001", b"11000000011001110000101000111101"), -- -1.04 + -2.57 = -3.61
	(b"11000000001100101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111111110000101000111101100", b"11000000100101110101110000101001"), -- -2.79 + -1.94 = -4.73
	(b"00111111101000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"00111111100111000010100011110110"), -- 1.27 + -0.05 = 1.22
	(b"00111111110001010001111010111000", b"00000000000000000000000000000000"),
	(b"01000000010111100001010001111011", b"01000000101000000101000111101100"), -- 1.54 + 3.47 = 5.01
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111010000000000000000000000", b"00111111000111000010100011110110"), -- -0.14 + 0.75 = 0.61
	(b"10111111010111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111001100001010001111010111", b"10111110001110000101000111101100"), -- -0.87 + 0.69 = -0.18
	(b"11000000000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011111010111000010100100", b"00111111111101000111101011100010"), -- -2.05 + 3.96 = 1.91
	(b"10111111010111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111111110101110000101001000", b"00111111100011001100110011001101"), -- -0.86 + 1.96 = 1.1
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001001011100001010001111", b"11000000101011111010111000010100"), -- -2.9 + -2.59 = -5.49
	(b"01000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000000011100001010001111011", b"00111111000101110000101000111100"), -- 2.81 + -2.22 = 0.59
	(b"11000000001011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111111101100001010001111010111", b"10111111101011100001010001111011"), -- -2.74 + 1.38 = -1.36
	(b"11000000001000111101011100001010", b"00000000000000000000000000000000"),
	(b"00111110110001111010111000010100", b"11000000000010101110000101001000"), -- -2.56 + 0.39 = -2.17
	(b"11000000000110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111100101011100001010001111", b"11000000011001011100001010010000"), -- -2.42 + -1.17 = -3.59
	(b"00111111001010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111111011100001010001111011", b"01000000001000010100011110101110"), -- 0.66 + 1.86 = 2.52
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000100100000000000000000000"), -- -1.2 + -3.3 = -4.5
	(b"00111111111011110101110000101001", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"00111111111101110000101000111101"), -- 1.87 + 0.06 = 1.93
	(b"01000000001111010111000010100100", b"00000000000000000000000000000000"),
	(b"01000000000100001010001111010111", b"01000000101001110000101000111110"), -- 2.96 + 2.26 = 5.22
	(b"10111110111010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000001100001010001111010111", b"11000000010011100001010001111011"), -- -0.46 + -2.76 = -3.22
	(b"01000000000111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111011100001010001111010111", b"00111111110001010001111010111000"), -- 2.48 + -0.94 = 1.54
	(b"00111110101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000000000110011001100110011"), -- 0.35 + 1.7 = 2.05
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111000110011001100110011000"), -- -2.6 + 2 = -0.6
	(b"01000000001101110000101000111101", b"00000000000000000000000000000000"),
	(b"11000000010011110101110000101001", b"10111110110000101000111101100000"), -- 2.86 + -3.24 = -0.38
	(b"00111111001111010111000010100100", b"00000000000000000000000000000000"),
	(b"10111111000101000111101011100001", b"00111110001000111101011100001100"), -- 0.74 + -0.58 = 0.16
	(b"00111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"01000000000000110011001100110011", b"01000000001111100001010001111011"), -- 0.92 + 2.05 = 2.97
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001001100110011001100110", b"11000000010100000000000000000000"), -- -2.6 + -0.65 = -3.25
	(b"00111111111000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111110111000010100011110110", b"00111101010011001100110011000000"), -- 1.77 + -1.72 = 0.05
	(b"11000000010000011110101110000101", b"00000000000000000000000000000000"),
	(b"10111111000011001100110011001101", b"11000000011001010001111010111000"), -- -3.03 + -0.55 = -3.58
	(b"01000000010101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"00111111111110000101000111101011"), -- 3.34 + -1.4 = 1.94
	(b"11000000001010000101000111101100", b"00000000000000000000000000000000"),
	(b"10111111101010100011110101110001", b"11000000011111010111000010100100"), -- -2.63 + -1.33 = -3.96
	(b"11000000010111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111111000010100011110101110", b"10111111110111000010100011110110"), -- -3.48 + 1.76 = -1.72
	(b"10111111101000101000111101011100", b"00000000000000000000000000000000"),
	(b"11000000010100010100011110101110", b"11000000100100010100011110101110"), -- -1.27 + -3.27 = -4.54
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110111000010100011111", b"10111111010001010001111010111000"), -- -3.2 + 2.43 = -0.77
	(b"01000000001110001111010111000011", b"00000000000000000000000000000000"),
	(b"10111111100101000111101011100001", b"00111111110111010111000010100101"), -- 2.89 + -1.16 = 1.73
	(b"01000000000111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111101000000000000000000000", b"01000000011011101011100001010010"), -- 2.48 + 1.25 = 3.73
	(b"00111111110110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111101010100011110101110001", b"00111110110000101000111101011100"), -- 1.71 + -1.33 = 0.38
	(b"01000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"00111101011101011100001010001111", b"01000000001001000111101011100001"), -- 2.51 + 0.06 = 2.57
	(b"11000000001000011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000000111010111000010100100", b"11000000100111111010111000010100"), -- -2.53 + -2.46 = -4.99
	(b"10111111110001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000101000111101011100", b"11000000001001000111101011100001"), -- -1.55 + -1.02 = -2.57
	(b"11000000010101011100001010001111", b"00000000000000000000000000000000"),
	(b"01000000001010011001100110011010", b"10111111001100001010001111010100"), -- -3.34 + 2.65 = -0.69
	(b"10111100001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110111001100110011001100110", b"10111110111010111000010100011110"), -- -0.01 + -0.45 = -0.46
	(b"01000000001000101000111101011100", b"00000000000000000000000000000000"),
	(b"10111111001100001010001111010111", b"00111111111011001100110011001100"), -- 2.54 + -0.69 = 1.85
	(b"11000000000000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000011110101110000101001000", b"00111111111011100001010001111100"), -- -2.06 + 3.92 = 1.86
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"10111111011000111101011100001010", b"10111110001000111101011100001000"), -- 0.73 + -0.89 = -0.16
	(b"11000000011011010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000010011010111000010100100"), -- -3.71 + 0.5 = -3.21
	(b"10111111111001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000011011000010100011110110", b"00111111111100001010001111011000"), -- -1.81 + 3.69 = 1.88
	(b"11000000011101010001111010111000", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"11000000011101111010111000010100"), -- -3.83 + -0.04 = -3.87
	(b"11000000010111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111000101000111101011100", b"11000000101001110000101000111110"), -- -3.45 + -1.77 = -5.22
	(b"10111111100001010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000000110001111010111000011", b"11000000010110111000010100011111"), -- -1.04 + -2.39 = -3.43
	(b"11000000011010000101000111101100", b"00000000000000000000000000000000"),
	(b"01000000000110001111010111000011", b"10111111100111101011100001010010"), -- -3.63 + 2.39 = -1.24
	(b"11000000011000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100101000111101011100", b"11000000110110101110000101001000"), -- -3.55 + -3.29 = -6.84
	(b"01000000011000011110101110000101", b"00000000000000000000000000000000"),
	(b"00111110111010111000010100011111", b"01000000011111110101110000101001"), -- 3.53 + 0.46 = 3.99
	(b"00111111101011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000010101000111101011100001", b"01000000100101011100001010001111"), -- 1.36 + 3.32 = 4.68
	(b"11000000001000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000010000010100011110101110", b"00111110111010111000010100100000"), -- -2.56 + 3.02 = 0.46
	(b"10111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000001111110101110000101001", b"11000000011100010100011110101110"), -- -0.78 + -2.99 = -3.77
	(b"01000000001111100001010001111011", b"00000000000000000000000000000000"),
	(b"00111110101100110011001100110011", b"01000000010101000111101011100001"), -- 2.97 + 0.35 = 3.32
	(b"10111111101110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000001111101011100001010010", b"11000000100011010111000010100100"), -- -1.44 + -2.98 = -4.42
	(b"01000000010000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001100111101011100001010", b"01000000101110111101011100001010"), -- 3.06 + 2.81 = 5.87
	(b"00111111010010100011110101110001", b"00000000000000000000000000000000"),
	(b"10111111010101000111101011100001", b"10111101001000111101011100000000"), -- 0.79 + -0.83 = -0.04
	(b"01000000001011010111000010100100", b"00000000000000000000000000000000"),
	(b"00111111111001111010111000010100", b"01000000100100001010001111010111"), -- 2.71 + 1.81 = 4.52
	(b"00111111000101110000101000111101", b"00000000000000000000000000000000"),
	(b"01000000000100111101011100001010", b"01000000001110011001100110011001"), -- 0.59 + 2.31 = 2.9
	(b"00111111010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101001000111101011100001010", b"00111111011000111101011100001011"), -- 0.85 + 0.04 = 0.89
	(b"00111111111000101000111101011100", b"00000000000000000000000000000000"),
	(b"00111111010000000000000000000000", b"01000000001000010100011110101110"), -- 1.77 + 0.75 = 2.52
	(b"10111111100111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111110110101110000101000111110"), -- -1.22 + 0.8 = -0.42
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101010011001100110011001101", b"01000000000111001100110011001101"), -- 2.5 + -0.05 = 2.45
	(b"10111110000011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000010100001010001111010111", b"11000000010110011001100110011010"), -- -0.14 + -3.26 = -3.4
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000001011001100110011001101"), -- -2.2 + -0.5 = -2.7
	(b"11000000000000001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000101110011110101110000101"), -- -2.01 + -3.8 = -5.81
	(b"10111110001000111101011100001010", b"00000000000000000000000000000000"),
	(b"10111110100010100011110101110001", b"10111110110111000010100011110110"), -- -0.16 + -0.27 = -0.43
	(b"11000000001010001111010111000011", b"00000000000000000000000000000000"),
	(b"01000000001101011100001010001111", b"00111110010011001100110011000000"), -- -2.64 + 2.84 = 0.2
	(b"00111110101000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000000000101000111101011100", b"01000000000101110000101000111101"), -- 0.32 + 2.04 = 2.36
	(b"01000000010001111010111000010100", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000000110101110000101000111"), -- 3.12 + -0.7 = 2.42
	(b"01000000011011101011100001010010", b"00000000000000000000000000000000"),
	(b"01000000010110001111010111000011", b"01000000111000111101011100001010"), -- 3.73 + 3.39 = 7.12
	(b"01000000010111101011100001010010", b"00000000000000000000000000000000"),
	(b"00111111001001100110011001100110", b"01000000100001000010100011110110"), -- 3.48 + 0.65 = 4.13
	(b"11000000011001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000010100010100011110101110", b"10111110101100110011001100110000"), -- -3.62 + 3.27 = -0.35
	(b"11000000000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000001000111101011100001", b"11000000100100001010001111010111"), -- -2.45 + -2.07 = -4.52
	(b"00111111111101011100001010001111", b"00000000000000000000000000000000"),
	(b"10111111100001111010111000010100", b"00111111010111000010100011110110"), -- 1.92 + -1.06 = 0.86
	(b"11000000001100111101011100001010", b"00000000000000000000000000000000"),
	(b"00111111010010100011110101110001", b"11000000000000010100011110101110"), -- -2.81 + 0.79 = -2.02
	(b"10111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"11000000011011101011100001010010", b"11000000011111001100110011001101"), -- -0.22 + -3.73 = -3.95
	(b"11000000011100001010001111010111", b"00000000000000000000000000000000"),
	(b"10111111110001100110011001100110", b"11000000101010011110101110000101"), -- -3.76 + -1.55 = -5.31
	(b"00111111111110000101000111101100", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111111110100011110101110000110"), -- 1.94 + -0.3 = 1.64
	(b"10111101010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110000101000111101100", b"01000000000101010001111010111001"), -- -0.05 + 2.38 = 2.33
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100101000111101011100", b"01000000100000101110000101001000"), -- 1.3 + 2.79 = 4.09
	(b"10111111101010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111111000000101000111101011100", b"10111111111011001100110011001101"), -- -1.34 + -0.51 = -1.85
	(b"11000000000010111000010100011111", b"00000000000000000000000000000000"),
	(b"10111101001000111101011100001010", b"11000000000011100001010001111011"), -- -2.18 + -0.04 = -2.22
	(b"00111111101000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000111101011100001010", b"01000000000100011110101110000101"), -- 1.25 + 1.03 = 2.28
	(b"01000000001001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111100001111010111000010100", b"00111111110000101000111101011100"), -- 2.58 + -1.06 = 1.52
	(b"10111111101101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111110100101000111101011100001", b"10111111100011110101110000101001"), -- -1.41 + 0.29 = -1.12
	(b"00111111010001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000011111010111000010100100", b"01000000100101111010111000010100"), -- 0.78 + 3.96 = 4.74
	(b"10111111001011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000011010111000010100011111", b"01000000010000000000000000000000"), -- -0.68 + 3.68 = 3
	(b"01000000000011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000000110111000010100011111", b"01000000100101010111000010100100"), -- 2.24 + 2.43 = 4.67
	(b"11000000000110100011110101110001", b"00000000000000000000000000000000"),
	(b"00111111011101011100001010001111", b"10111111101110011001100110011010"), -- -2.41 + 0.96 = -1.45
	(b"01000000001010001111010111000011", b"00000000000000000000000000000000"),
	(b"00111111011100001010001111010111", b"01000000011001010001111010111001"), -- 2.64 + 0.94 = 3.58
	(b"01000000001111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011100001010001111011", b"10111111010001010001111010111000"), -- 2.95 + -3.72 = -0.77
	(b"01000000000011100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000001100101000111101011100", b"01000000101000000101000111101100"), -- 2.22 + 2.79 = 5.01
	(b"10111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000100110111000010100011110"), -- -1.56 + -3.3 = -4.86
	(b"00111111101000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111110011001100110011010", b"10111111001100110011001100110100"), -- 1.25 + -1.95 = -0.7
	(b"00111111101000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"00111111010111101011100001010010"), -- 1.25 + -0.38 = 0.87
	(b"10111111111011100001010001111011", b"00000000000000000000000000000000"),
	(b"11000000000111001100110011001101", b"11000000100010011110101110000101"), -- -1.86 + -2.45 = -4.31
	(b"10111111011010111000010100011111", b"00000000000000000000000000000000"),
	(b"11000000000010001111010111000011", b"11000000010000111101011100001011"), -- -0.92 + -2.14 = -3.06
	(b"00111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"10111111010101110000101000111101", b"10111111000011110101110000101000"), -- 0.28 + -0.84 = -0.56
	(b"01000000010111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110101110000101000111101100", b"01000000010001011100001010010000"), -- 3.45 + -0.36 = 3.09
	(b"00111111100110000101000111101100", b"00000000000000000000000000000000"),
	(b"11000000011101000111101011100001", b"11000000001010000101000111101011"), -- 1.19 + -3.82 = -2.63
	(b"10111111111111101011100001010010", b"00000000000000000000000000000000"),
	(b"10111111001110101110000101001000", b"11000000001011100001010001111011"), -- -1.99 + -0.73 = -2.72
	(b"01000000000101110000101000111101", b"00000000000000000000000000000000"),
	(b"10111111001101011100001010001111", b"00111111110100110011001100110010"), -- 2.36 + -0.71 = 1.65
	(b"01000000010111000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000001100011110101110000101", b"01000000110001110000101000111110"), -- 3.44 + 2.78 = 6.22
	(b"11000000001101010001111010111000", b"00000000000000000000000000000000"),
	(b"11000000011101010001111010111000", b"11000000110101010001111010111000"), -- -2.83 + -3.83 = -6.66
	(b"01000000000111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110101110000101001000", b"00111111100111101011100001010010"), -- 2.45 + -1.21 = 1.24
	(b"01000000011100010100011110101110", b"00000000000000000000000000000000"),
	(b"10111110110000101000111101011100", b"01000000010110001111010111000010"), -- 3.77 + -0.38 = 3.39
	(b"11000000000100101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000010000110011001100110011", b"00111111010000101000111101011100"), -- -2.29 + 3.05 = 0.76
	(b"11000000011111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111101100011110101110000101001", b"11000000011101111010111000010101"), -- -3.94 + 0.07 = -3.87
	(b"01000000001100001010001111010111", b"00000000000000000000000000000000"),
	(b"11000000010111000010100011110110", b"10111111001011100001010001111100"), -- 2.76 + -3.44 = -0.68
	(b"00111111111100011110101110000101", b"00000000000000000000000000000000"),
	(b"11000000000011100001010001111011", b"10111110101010001111010111000100"), -- 1.89 + -2.22 = -0.33
	(b"01000000001000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111110111010111000010100100", b"01000000100010000000000000000000"), -- 2.52 + 1.73 = 4.25
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000001111100001010001111011", b"01000000010101100110011001100110"), -- 0.38 + 2.97 = 3.35
	(b"11000000010010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111011100001010001111011", b"11000000101000000101000111101100"), -- -3.15 + -1.86 = -5.01
	(b"00111111101100011110101110000101", b"00000000000000000000000000000000"),
	(b"00111111001010001111010111000011", b"01000000000000110011001100110011"), -- 1.39 + 0.66 = 2.05
	(b"01000000000111100001010001111011", b"00000000000000000000000000000000"),
	(b"01000000001100011110101110000101", b"01000000101010000000000000000000"), -- 2.47 + 2.78 = 5.25
	(b"10111110100011110101110000101001", b"00000000000000000000000000000000"),
	(b"11000000010100111101011100001010", b"11000000011001011100001010001111"), -- -0.28 + -3.31 = -3.59
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000010110011001100110011010"), -- 1.7 + 1.7 = 3.4
	(b"01000000011001010001111010111000", b"00000000000000000000000000000000"),
	(b"10111111010001010001111010111000", b"01000000001100111101011100001010"), -- 3.58 + -0.77 = 2.81
	(b"00111111001110101110000101001000", b"00000000000000000000000000000000"),
	(b"11000000001111000010100011110110", b"11000000000011010111000010100100"), -- 0.73 + -2.94 = -2.21
	(b"01000000011111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100101000111101011100", b"00111111100101000111101011100010"), -- 3.95 + -2.79 = 1.16
	(b"01000000001000001010001111010111", b"00000000000000000000000000000000"),
	(b"10111101111101011100001010001111", b"01000000000110001111010111000011"), -- 2.51 + -0.12 = 2.39
	(b"00111110110000101000111101011100", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011010111000010100011110"), -- 0.38 + 3.3 = 3.68
	(b"00111111001110000101000111101100", b"00000000000000000000000000000000"),
	(b"00111111100111010111000010100100", b"00111111111110011001100110011010"), -- 0.72 + 1.23 = 1.95
	(b"11000000010001011100001010001111", b"00000000000000000000000000000000"),
	(b"00111111100100110011001100110011", b"10111111111110000101000111101011"), -- -3.09 + 1.15 = -1.94
	(b"00111111101111000010100011110110", b"00000000000000000000000000000000"),
	(b"00111111011111010111000010100100", b"01000000000111010111000010100100"), -- 1.47 + 0.99 = 2.46
	(b"11000000010000111101011100001010", b"00000000000000000000000000000000"),
	(b"11000000001101111010111000010100", b"11000000101111011100001010001111"), -- -3.06 + -2.87 = -5.93
	(b"00111111011000111101011100001010", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000011001011100001010010000"), -- 0.89 + 2.7 = 3.59
	(b"00111111010100011110101110000101", b"00000000000000000000000000000000"),
	(b"10111110101010001111010111000011", b"00111110111110101110000101000111"), -- 0.82 + -0.33 = 0.49
	(b"10111110011000010100011110101110", b"00000000000000000000000000000000"),
	(b"00111111100111010111000010100100", b"00111111100000010100011110101110"), -- -0.22 + 1.23 = 1.01
	(b"00111111010011110101110000101001", b"00000000000000000000000000000000"),
	(b"01000000001011000010100011110110", b"01000000011000000000000000000000"), -- 0.81 + 2.69 = 3.5
	(b"10111110101111010111000010100100", b"00000000000000000000000000000000"),
	(b"11000000001000011110101110000101", b"11000000001110011001100110011010"), -- -0.37 + -2.53 = -2.9
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001110000101000111101", b"01000000101101101011100001010010"), -- 2.1 + 3.61 = 5.71
	(b"11000000010011000010100011110110", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000100011111010111000010100"), -- -3.19 + -1.3 = -4.49
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001000111101011100001", b"11000000011111100001010001111010"), -- -1.4 + -2.57 = -3.97
	(b"11000000001011000010100011110110", b"00000000000000000000000000000000"),
	(b"01000000011000111101011100001010", b"00111111010111101011100001010000"), -- -2.69 + 3.56 = 0.87
	(b"11000000001101000111101011100001", b"00000000000000000000000000000000"),
	(b"00111111101101000111101011100001", b"10111111101101000111101011100001"), -- -2.82 + 1.41 = -1.41
	(b"10111111110001111010111000010100", b"00000000000000000000000000000000"),
	(b"01000000001111101011100001010010", b"00111111101101011100001010010000"), -- -1.56 + 2.98 = 1.42
	(b"00111111100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000111000010100011110110", b"01000000011001011100001010010000"), -- 1.15 + 2.44 = 3.59
	(b"00111111100001111010111000010100", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000000101110000101000111101"), -- 1.06 + 1.3 = 2.36
	(b"00111111110010001111010111000011", b"00000000000000000000000000000000"),
	(b"11000000001011110101110000101001", b"10111111100101011100001010001111"), -- 1.57 + -2.74 = -1.17

	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- -0 + 1.7 = 1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- 0 + 0.4 = 0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- 0 + 0.7 = 0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- 0 + -2.8 = -2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- 0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- 0 + -0.2 = -0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- -0 + 3.6 = 3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- 0 + 2.7 = 2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- -0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- -0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- -0 + 3.3 = 3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- -0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- -0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- 0 + -1.7 = -1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- -0 + -2.3 = -2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- -0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- 0 + -1.7 = -1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- 0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- 0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- 0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- 0 + 0.8 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- 0 + -2.8 = -2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- -0 + 2.9 = 2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- -0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- -0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- 0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- 0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- 0 + 0.2 = 0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- -0 + -2.5 = -2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- 0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- -0 + 0.4 = 0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- -0 + -2.3 = -2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- 0 + -2.7 = -2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- -0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- -0 + 1.2 = 1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- -0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- -0 + 0.3 = 0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- 0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- -0 + -2.7 = -2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- 0 + -2.7 = -2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- -0 + -1.2 = -1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- -0 + 1 = 1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- -0 + 1.1 = 1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- 0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- -0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- -0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- 0 + 0.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- 0 + -3.1 = -3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- -0 + 1 = 1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- 0 + 0.4 = 0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- -0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- 0 + 0.4 = 0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- -0 + -2.5 = -2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- 0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- -0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- 0 + -1.9 = -1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- 0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- 0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- -0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- -0 + 0.5 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- 0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010110011001100110011010"), -- 0 + -3.4 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- 0 + 0.9 = 0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- -0 + 0.1 = 0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- -0 + 1 = 1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- 0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010110011001100110011010"), -- -0 + -3.4 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- -0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- 0 + 1 = 1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- -0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- 0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- 0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- -0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- -0 + -0.2 = -0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- -0 + -1.2 = -1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- -0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- 0 + 2.7 = 2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- 0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- -0 + 0.7 = 0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- -0 + 0.1 = 0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- -0 + -2.5 = -2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- -0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- -0 + -1.8 = -1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- 0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- -0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- 0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- 0 + 3.8 = 3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- 0 + -2.8 = -2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- -0 + -2 = -2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- -0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- 0 + 3.8 = 3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- -0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- 0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- -0 + -1.7 = -1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- -0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- 0 + 3.4 = 3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- 0 + 0.2 = 0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- -0 + -1.2 = -1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- 0 + -2.8 = -2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- 0 + -3.1 = -3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- -0 + 1.4 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- 0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- -0 + -1.8 = -1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- 0 + -3 = -3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- -0 + 3.7 = 3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- 0 + 3.6 = 3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- -0 + -3.3 = -3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- -0 + -3.3 = -3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- 0 + 2 = 2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- -0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- 0 + -1.7 = -1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- -0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- -0 + -2.8 = -2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- -0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- 0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- -0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- 0 + -2.7 = -2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- -0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- 0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- -0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- 0 + -1.2 = -1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- 0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- -0 + 0.5 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- 0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- -0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- -0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- 0 + -3 = -3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- -0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- 0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- 0 + -2.7 = -2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- -0 + 3.1 = 3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- 0 + 2.6 = 2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- -0 + -1.8 = -1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- 0 + 3.6 = 3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- -0 + 1.7 = 1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- -0 + -3.9 = -3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- 0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- 0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- -0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- 0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- -0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- -0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- -0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- -0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- 0 + 0.4 = 0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- -0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- 0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- -0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- 0 + 0.9 = 0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- -0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- 0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- -0 + 3.6 = 3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- -0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- -0 + 3.5 = 3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- 0 + 1 = 1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- -0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- -0 + 0.7 = 0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- -0 + -3.3 = -3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- 0 + -1.2 = -1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- 0 + 0.5 = 0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- -0 + 0.5 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- 0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- 0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- -0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- -0 + 0.7 = 0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- -0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- -0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- -0 + -3.7 = -3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- -0 + 0.7 = 0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- -0 + -0.3 = -0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- -0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- -0 + -2.3 = -2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- 0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- -0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- 0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- 0 + 1.5 = 1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- -0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- -0 + 0.7 = 0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- -0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- 0 + -1.6 = -1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- -0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- 0 + 0.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- 0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- -0 + 0.7 = 0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- 0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- -0 + -0.2 = -0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- -0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010110011001100110011010"), -- -0 + -3.4 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- -0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- -0 + -0.2 = -0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- -0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- -0 + 1.7 = 1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- -0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- -0 + -2.6 = -2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- 0 + 1.4 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- 0 + -1.8 = -1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- -0 + -0.2 = -0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- -0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- -0 + 3.5 = 3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- -0 + -2.8 = -2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- 0 + -1.9 = -1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- 0 + -2.8 = -2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- -0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- 0 + 3.2 = 3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- -0 + 0.3 = 0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- 0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- 0 + -1.9 = -1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- 0 + -3.6 = -3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- 0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- -0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- 0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010110011001100110011010"), -- 0 + -3.4 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- 0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- 0 + -1.6 = -1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- 0 + 3.6 = 3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- -0 + 0.5 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- 0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- 0 + 3.8 = 3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- -0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- -0 + 0.5 = 0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- -0 + -2.3 = -2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- -0 + 1.3 = 1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- -0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- -0 + 0.4 = 0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- -0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- 0 + -1.7 = -1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- -0 + 1.2 = 1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- -0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- -0 + 1.1 = 1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- -0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- -0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- 0 + 3.5 = 3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- 0 + 3.2 = 3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- 0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- -0 + 3.7 = 3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- 0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- -0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- -0 + 0.5 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- 0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- -0 + -1.9 = -1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- 0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- 0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- -0 + 0.1 = 0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- -0 + 2.3 = 2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- 0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- 0 + 2 = 2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- -0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- 0 + 1 = 1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- 0 + -1.8 = -1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- 0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- 0 + -2.7 = -2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- -0 + -1.8 = -1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- 0 + -1.6 = -1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- 0 + 2.7 = 2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111110110011001100110011010"), -- -0 + 1.7 = 1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- 0 + -3.2 = -3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- -0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- -0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- 0 + -3.6 = -3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- 0 + 3.2 = 3.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- 0 + 2.4 = 2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- 0 + -1.2 = -1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- 0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- 0 + -3.6 = -3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- -0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- -0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001011001100110011001101"), -- -0 + 2.7 = 2.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000001000000000000000000000"), -- -0 + 2.5 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- 0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10000000000000000000000000000000"), -- -0 + -0 = -0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- -0 + 1.1 = 1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- 0 + -1.7 = -1.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- 0 + -3.9 = -3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- -0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- 0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- 0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- -0 + -2.9 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- -0 + 2.1 = 2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- 0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- -0 + 3.7 = 3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- 0 + -3.2 = -3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- 0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- 0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- 0 + -2.1 = -2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- 0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- -0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- -0 + -3.6 = -3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- 0 + 1.4 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- 0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- 0 + 2.6 = 2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- 0 + -0.2 = -0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- -0 + 1.4 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- 0 + 0.5 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- -0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- 0 + -3 = -3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- -0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- 0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- -0 + 3.7 = 3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- 0 + 3.6 = 3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- -0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- 0 + -1 = -1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111110110011001100110011010"), -- -0 + -1.7 = -1.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- 0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- 0 + 0.7 = 0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- 0 + 2 = 2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- 0 + -3.5 = -3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- -0 + 0.8 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- -0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000000001100110011001100110"), -- -0 + -2.1 = -2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110010011001100110011001101"), -- -0 + -0.2 = -0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- -0 + 2.4 = 2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- -0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010100110011001100110011"), -- 0 + -3.3 = -3.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- -0 + 2.6 = 2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- -0 + -0.6 = -0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- 0 + -3.7 = -3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- -0 + 0.9 = 0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- -0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100110011001100110011010"), -- 0 + 1.2 = 1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- 0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011000000000000000000000"), -- -0 + -3.5 = -3.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- 0 + -2.7 = -2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- 0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- -0 + 1.4 = 1.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- -0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- 0 + -2 = -2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- -0 + 3.6 = 3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- -0 + 3.8 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- 0 + 0.2 = 0.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- -0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100000000000000000000000"), -- -0 + -1 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- -0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- -0 + 0 = 0
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011000000000000000000000"), -- -0 + 3.5 = 3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- 0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111000110011001100110011010"), -- 0 + -0.6 = -0.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- -0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- -0 + 3.4 = 3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- 0 + 2.1 = 2.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- -0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001011001100110011001101"), -- -0 + -2.7 = -2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- 0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- -0 + -3 = -3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001000000000000000000000"), -- 0 + -2.5 = -2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- 0 + 0.9 = 0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- 0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111110011001100110011001101"), -- 0 + -1.6 = -1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111101100110011001100110011"), -- -0 + 1.4 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111000110011001100110011010"), -- 0 + 0.6 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001001100110011001100110"), -- 0 + -2.6 = -2.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- -0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- -0 + 1.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- 0 + 1 = 1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010100110011001100110011"), -- 0 + 3.3 = 3.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000011011001100110011001101"), -- -0 + -3.7 = -3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011110011001100110011010"), -- -0 + 3.9 = 3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- 0 + 1.8 = 1.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111011001100110011001100110"), -- -0 + 0.9 = 0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011110011001100110011010"), -- -0 + -3.9 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- 0 + 0.7 = 0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- -0 + -1.2 = -1.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- -0 + -2 = -2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- -0 + -3.1 = -3.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111111100110011001100110011"), -- 0 + -1.9 = -1.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111110011001100110011001101"), -- -0 + 1.6 = 1.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000000000000000000000000"), -- -0 + -2 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000011100110011001100110011"), -- -0 + 3.8 = 3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- -0 + 2.8 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- 0 + 3.6 = 3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111110110011001100110011001101"), -- 0 + 0.4 = 0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110100110011001100110011010"), -- -0 + 0.3 = 0.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- -0 + 2.9 = 2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- -0 + -2.8 = -2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111111001100110011001100110"), -- -0 + -1.8 = -1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111100011001100110011001101"), -- 0 + 1.1 = 1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- -0 + -3.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- -0 + -2.4 = -2.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000001110011001100110011010"), -- -0 + 2.9 = 2.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000001100110011001100110011"), -- 0 + 2.8 = 2.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010011001100110011001101"), -- -0 + -3.2 = -3.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011001100110011001100110"), -- 0 + 3.6 = 3.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- -0 + -0.8 = -0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111001100110011001100110"), -- -0 + 1.8 = 1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- 0 + -0.7 = -0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111110010011001100110011001101"), -- -0 + 0.2 = 0.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- -0 + -0.1 = -0.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- -0 + -0.4 = -0.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- 0 + 0.7 = 0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100011001100110011001101"), -- 0 + -1.1 = -1.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111001100110011001100110011"), -- -0 + -0.7 = -0.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- -0 + 1.5 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100000000000000000000000"), -- 0 + 1 = 1

	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000101001100110011001100110"), -- 3.1 + 2.1 = 5.2
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000101011001100110011001101"), -- -2.4 + -3 = -5.4
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000000110011001100110011001"), -- 2.3 + 0.1 = 2.4
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"10111110110011001100110011001000"), -- -2.1 + 1.7 = -0.4
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000100100000000000000000000"), -- -0.6 + -3.9 = -4.5
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000100000000000000000000000"), -- 1.2 + 2.8 = 4
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000010011001100110011001101"), -- -2.8 + -0.4 = -3.2
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111001100110011001100110100"), -- -2.2 + 1.5 = -0.7
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111111100000000000000000000000"), -- -1.4 + 0.4 = -1
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000101111001100110011001100"), -- -2.1 + -3.8 = -5.9
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000011110011001100110011010"), -- -3.3 + -0.6 = -3.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010110011001100110011010"), -- 0 + 3.4 = 3.4
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000100001100110011001100110"), -- 3.6 + 0.6 = 4.2
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001110011001100110011001"), -- 0.3 + 2.6 = 2.9
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"), -- -3.2 + 3.2 = 0
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111001100110011001100110011"), -- -0.8 + 1.5 = 0.7
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000101011001100110011001101"), -- 1.5 + 3.9 = 5.4
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000100001100110011001100110"), -- 2.8 + 1.4 = 4.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"00111110010011001100110011010000"), -- 3.2 + -3 = 0.2
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000000000000000000000000000"), -- -1.3 + 3.3 = 2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111000000000000000000000001"), -- 0.7 + -1.2 = -0.5
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000000000000000000000000000"), -- -1.8 + -0.2 = -2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000001001100110011001100110"), -- 2 + 0.6 = 2.6
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000111000000000000000000000"), -- 3.9 + 3.1 = 7
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000010110011001100110011001"), -- 3.6 + -0.2 = 3.4
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000101001100110011001100110"), -- -3.9 + -1.3 = -5.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"00111111110000000000000000000000"), -- 2.8 + -1.3 = 1.5
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000101111001100110011001101"), -- 3 + 2.9 = 5.9
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"00111110110011001100110011001100"), -- 1.9 + -1.5 = 0.4
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000100000110011001100110011"), -- 0.7 + 3.4 = 4.1
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010100110011001100110011"), -- -0.2 + -3.1 = -3.3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111110110011001100110011001110"), -- 0.7 + -1.1 = -0.4
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"00111111111001100110011001100110"), -- 3.1 + -1.3 = 1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000110011001100110011010"), -- 0 + 2.4 = 2.4
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000000001100110011001100110"), -- -0.9 + 3 = 2.1
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000111101100110011001100110"), -- 3.9 + 3.8 = 7.7
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000010011001100110011001100"), -- 0.4 + -3.6 = -3.2
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000010110011001100110011010"), -- -3 + -0.4 = -3.4
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000110001100110011001100110"), -- 2.4 + 3.8 = 6.2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111011001100110011001100110"), -- 0.2 + 0.7 = 0.9
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110011001100110011001101"), -- 0.1 + 1.5 = 1.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000001001100110011001100110"), -- 2 + 0.6 = 2.6
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000001100110011001100110011"), -- -2.8 + -0 = -2.8
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000001001100110011001100110"), -- 3.2 + -0.6 = 2.6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000001000000000000000000000"), -- 0.8 + -3.3 = -2.5
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111111110110011001100110011010"), -- -2 + 0.3 = -1.7
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000010011001100110011001101"), -- 1.7 + 1.5 = 3.2
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010011001100110011001100"), -- 0.1 + 3.1 = 3.2
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111110110011001100110011010"), -- -1.6 + -0.1 = -1.7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000011110011001100110011010"), -- 3.7 + 0.2 = 3.9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000101000000000000000000000"), -- 2.9 + 2.1 = 5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000011110011001100110011010"), -- -0.7 + -3.2 = -3.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000001001100110011001100110"), -- 3 + -0.4 = 2.6
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111111000110011001100110011000"), -- -3.1 + 2.5 = -0.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111101001100110011001100110"), -- -1.3 + 2.6 = 1.3
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000011011001100110011001101"), -- 0.3 + 3.4 = 3.7
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000000100110011001100110100"), -- 0.6 + -2.9 = -2.3
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000110000000000000000000000"), -- -3.2 + -2.8 = -6
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"), -- -3 + 3 = 0
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000111100000000000000000000"), -- -3.9 + -3.6 = -7.5
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111110000000000000000000000"), -- 1 + 0.5 = 1.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000110100110011001100110011"), -- 3.5 + 3.1 = 6.6
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000101111001100110011001100"), -- -3.6 + -2.3 = -5.9
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100110011001100110011010"), -- 1.3 + 3.5 = 4.8
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111001100110011001100110100"), -- 2.6 + -3.3 = -0.7
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000011001100110011001100110"), -- -1.5 + -2.1 = -3.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111111110110011001100110011010"), -- -2 + 0.3 = -1.7
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000001000000000000000000000"), -- -1 + -1.5 = -2.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000100001100110011001100110"), -- 2.5 + 1.7 = 4.2
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111101001100110011001100110"), -- -1.5 + 2.8 = 1.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000001100110011001100110100"), -- 0.6 + 2.2 = 2.8
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000100001100110011001100110"), -- 1.2 + 3 = 4.2
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000111010011001100110011010"), -- -3.6 + -3.7 = -7.3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000101100110011001100110011"), -- -2.5 + -3.1 = -5.6
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00111111011001100110011001100110"), -- -1.6 + 2.5 = 0.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111010011001100110011001100"), -- 3 + -3.8 = -0.8
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000110011001100110011001101"), -- -2.5 + -3.9 = -6.4
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000110101100110011001100110"), -- 3.2 + 3.5 = 6.7
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111010011001100110011001101"), -- 0.2 + 0.6 = 0.8
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000111000000000000000000000"), -- -3.2 + -3.8 = -7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000010110011001100110011010"), -- 3.4 + -0 = 3.4
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111111111001100110011001100111"), -- -2.7 + 0.9 = -1.8
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101010011001100110011010"), -- 2.8 + 2.5 = 5.3
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000101110011001100110011010"), -- -3.1 + -2.7 = -5.8
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111111100011001100110011001100"), -- 2.3 + -1.2 = 1.1
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111010011001100110011001100"), -- 1.1 + -1.9 = -0.8
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111110100110011001100110011000"), -- 1.6 + -1.9 = -0.3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"10111110110011001100110011001101"), -- -0.5 + 0.1 = -0.4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000110110011001100110011010"), -- -3.8 + -3 = -6.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"00111110010011001100110011010000"), -- 3.7 + -3.5 = 0.2
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111110011001100110011001101"), -- 2.2 + -0.6 = 1.6
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000100100000000000000000000"), -- -2.9 + -1.6 = -4.5
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111111100000000000000000000000"), -- 1.7 + -0.7 = 1
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111111101100110011001100110010"), -- 1.7 + -3.1 = -1.4
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000000011100110011001100110011"), -- 3.3 + 0.5 = 3.8
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111101100110011001100110010"), -- 1.2 + -2.6 = -1.4
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000001001100110011001100110"), -- -1.2 + 3.8 = 2.6
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010000000000000000000000"), -- -0.3 + 3.3 = 3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000001110011001100110011010"), -- -0.6 + -2.3 = -2.9
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000011001100110011001100110"), -- 3.6 + -0 = 3.6
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000010110011001100110011010"), -- -1 + -2.4 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000010001100110011001100110"), -- 0 + 3.1 = 3.1
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"00111111110000000000000000000000"), -- -1.7 + 3.2 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010001100110011001100110"), -- 0 + -3.1 = -3.1
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111010011001100110011010000"), -- 3.1 + -3.9 = -0.8
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111000000000000000000000000"), -- -1 + 1.5 = 0.5
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000101000000000000000000000"), -- -2.9 + -2.1 = -5
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111110010011001100110011001110"), -- -0.4 + 0.6 = 0.2
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000010000000000000000000000"), -- -2.7 + -0.3 = -3
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111100000000000000000000000"), -- -2.9 + 3.9 = 1
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101111001100110011001100"), -- -3.3 + -2.6 = -5.9
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000010011001100110011001101"), -- 2 + 1.2 = 3.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"00111111000000000000000000000000"), -- 2.8 + -2.3 = 0.5
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000001100110011001100110100"), -- 1.1 + 1.7 = 2.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111100000000000000000000000"), -- 3.7 + -2.7 = 1
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000110001100110011001100110"), -- 3 + 3.2 = 6.2
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000100000000000000000000000"), -- -3 + -1 = -4
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00111110100110011001100110011000"), -- -2.8 + 3.1 = 0.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111011001100110011001100111"), -- 0.6 + 0.3 = 0.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000001011001100110011001101"), -- -0.3 + -2.4 = -2.7
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000001110011001100110011010"), -- -0.7 + -2.2 = -2.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000110101100110011001100110"), -- 2.8 + 3.9 = 6.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111110110011001100110011001000"), -- 2.2 + -2.6 = -0.4
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111011001100110011001100110"), -- -2.8 + 1.9 = -0.9
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111101110011001100110011000000"), -- 2.6 + -2.5 = 0.0999999
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111100000000000000000000000"), -- 1 + -0 = 1
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111110100110011001100110011100"), -- 2.2 + -1.9 = 0.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000110000000000000000000000"), -- -3.6 + -2.4 = -6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"00111111100011001100110011001100"), -- 3.3 + -2.2 = 1.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000011001100110011001101"), -- 0 + 2.2 = 2.2
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111111010011001100110011001110"), -- -1.9 + 2.7 = 0.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111101100110011001100110100"), -- -0.3 + 1.7 = 1.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000010000000000000000000000"), -- -1.1 + -1.9 = -3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000001100110011001100110011"), -- 0.9 + 1.9 = 2.8
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000101110011001100110011010"), -- -2.9 + -2.9 = -5.8
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000100001100110011001100110"), -- -3.5 + -0.7 = -4.2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111011001100110011001100110"), -- -2.5 + 1.6 = -0.9
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111110100110011001100110100000"), -- -2.6 + 2.9 = 0.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111101001100110011001101000"), -- 2.1 + -3.4 = -1.3
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000001011001100110011001101"), -- -1.1 + -1.6 = -2.7
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000011001100110011001100111"), -- 2.9 + 0.7 = 3.6
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000000011001100110011001101"), -- 1.6 + 0.6 = 2.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101001100110011001100110"), -- 0 + -1.3 = -1.3
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000101011001100110011001100"), -- 3.1 + 2.3 = 5.4
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"), -- -3.1 + 3.1 = 0
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111110100110011001100110011000"), -- -1.8 + 1.5 = -0.3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"10111110100110011001100110011000"), -- -2.5 + 2.2 = -0.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101010011001100110011010"), -- 2.8 + 2.5 = 5.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000110101100110011001100110"), -- 3.4 + 3.3 = 6.7
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"11000000001001100110011001100110"), -- -2.5 + -0.1 = -2.6
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111101001100110011001100110"), -- 1.4 + -0.1 = 1.3
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111111110110011001100110011010"), -- 1 + -2.7 = -1.7
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"00111111100000000000000000000000"), -- 3.3 + -2.3 = 1
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000000001100110011001100110"), -- -2.6 + 0.5 = -2.1
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000100001100110011001100110"), -- 2 + 2.2 = 4.2
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000010110011001100110011010"), -- -1 + -2.4 = -3.4
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111101110011001100110011000000"), -- -3.2 + 3.3 = 0.0999999
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00111111010011001100110011001100"), -- -1.7 + 2.5 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000011001100110011001100110"), -- -3.8 + 0.2 = -3.6
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000101011001100110011001101"), -- -3.7 + -1.7 = -5.4
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000011001100110011001100110"), -- -2.8 + -0.8 = -3.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111111111111111111111111111111"), -- -0.1 + 2.1 = 2
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111001100110011001100110010"), -- 2.6 + -1.9 = 0.7
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000011110011001100110011010"), -- -1.7 + -2.2 = -3.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000000011001100110011001101"), -- -0.3 + -1.9 = -2.2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000100101100110011001100110"), -- -1.1 + -3.6 = -4.7
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000100100110011001100110011"), -- 2.8 + 1.8 = 4.6
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"10111110100110011001100110100000"), -- -2.9 + 2.6 = -0.3
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110110011001100110011010"), -- 3.2 + 3.6 = 6.8
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111010011001100110011001100"), -- 1.9 + -1.1 = 0.8
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000000110011001100110011010"), -- -1.6 + -0.8 = -2.4
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000011001100110011001100110"), -- 1.3 + 2.3 = 3.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000001110011001100110011010"), -- 3.5 + -0.6 = 2.9
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111101100110011001100110100"), -- -3.4 + 2 = -1.4
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111010011001100110011001101"), -- 0.8 + -0 = 0.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"00111111100110011001100110011001"), -- 1.4 + -0.2 = 1.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000100001100110011001100110"), -- 2.8 + 1.4 = 4.2
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000000011001100110011001100"), -- -1.4 + 3.6 = 2.2
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000111000110011001100110100"), -- 3.7 + 3.4 = 7.1
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111110010011001100110011001101"), -- -0.4 + 0.2 = -0.2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111111010011001100110011001101"), -- 0.2 + 0.6 = 0.8
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000110101100110011001100110"), -- -3.2 + -3.5 = -6.7
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111111111100110011001100110011"), -- 1.8 + 0.1 = 1.9
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"10111101110011001100110011100000"), -- -3.4 + 3.3 = -0.1
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000100010011001100110011010"), -- -1.7 + -2.6 = -4.3
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111111001100110011001100110100"), -- 3 + -3.7 = -0.7
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111101001100110011001100110"), -- 3.8 + -2.5 = 1.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000001000000000000000000000"), -- -0.6 + -1.9 = -2.5
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111010011001100110011001100"), -- -3 + 3.8 = 0.8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000110000110011001100110011"), -- 3.6 + 2.5 = 6.1
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000100000000000000000000000"), -- -0.9 + -3.1 = -4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111110110011001100110011010000"), -- 3 + -3.4 = -0.4
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111100011001100110011001100"), -- -0.7 + 1.8 = 1.1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111000110011001100110011010"), -- 0.6 + -1.2 = -0.6
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000000010000000000000000000000"), -- 3.8 + -0.8 = 3
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111110110011001100110011001100"), -- 1.4 + -1 = 0.4
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111101110011001100110011001101"), -- 0.1 + -0.2 = -0.1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111110100110011001100110011000"), -- 2.5 + -2.8 = -0.3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111000000000000000000000000"), -- -0.5 + 1 = 0.5
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111110110011001100110011001"), -- 2.8 + -1.1 = 1.7
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111111111001100110011001100110"), -- 0.2 + -2 = -1.8
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000100101100110011001100110"), -- -1.3 + -3.4 = -4.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111110011001100110011001100"), -- 2.2 + -3.8 = -1.6
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111111001100110011001100110"), -- -0.3 + -1.5 = -1.8
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000100010011001100110011010"), -- -2.7 + -1.6 = -4.3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111000000000000000000000000"), -- 2.6 + -2.1 = 0.5
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111100011001100110011001101"), -- -0.5 + -0.6 = -1.1
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000001100110011001100110011"), -- -1 + 3.8 = 2.8
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000100100110011001100110100"), -- 2.4 + 2.2 = 4.6
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111111011001100110011001100100"), -- -1.2 + 2.1 = 0.9
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"00111111000000000000000000000000"), -- 2.2 + -1.7 = 0.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000000000000000000000000"), -- 0.4 + -2.4 = -2
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000000001100110011001100110"), -- 3.6 + -1.5 = 2.1
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000011001100110011001100111"), -- -3.9 + 0.3 = -3.6
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000101001100110011001100110"), -- -1.5 + -3.7 = -5.2
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111110010011001100110011001000"), -- -2.1 + 1.9 = -0.2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111111100110011001100110100"), -- -1.2 + -0.7 = -1.9
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111111000000000000000000000000"), -- -3.1 + 3.6 = 0.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101000000000000000000000"), -- 2.5 + 2.5 = 5
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000010110011001100110011010"), -- 1.7 + 1.7 = 3.4
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111111110011001100110011001100"), -- 1.9 + -0.3 = 1.6
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000110000000000000000000000"), -- -2.9 + -3.1 = -6
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000100011001100110011001101"), -- 2.4 + 2 = 4.4
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000100001100110011001100110"), -- 3.6 + 0.6 = 4.2
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000101011001100110011001101"), -- 2.7 + 2.7 = 5.4
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111001100110011001100110100"), -- -2.8 + 3.5 = 0.7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111110011001100110011001100"), -- -2.8 + 1.2 = -1.6
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000100100000000000000000000"), -- -0.8 + -3.7 = -4.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"10111111100011001100110011001110"), -- 2.1 + -3.2 = -1.1
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111001100110011001100110010"), -- -1.9 + 2.6 = 0.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111100110011001100110011010"), -- 2.2 + -1 = 1.2
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000110100110011001100110011"), -- -3.8 + -2.8 = -6.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001001100110011001100111"), -- -0.1 + 2.7 = 2.6
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111101110011001100110011000000"), -- 2.8 + -2.7 = 0.0999999
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111111001100110011001100110011"), -- 1.4 + -0.7 = 0.7
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"00111110010011001100110011010000"), -- -3 + 3.2 = 0.2
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111101110011001100110011100000"), -- 3.8 + -3.9 = -0.1
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000100100110011001100110011"), -- -3.5 + -1.1 = -4.6
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111110010011001100110011001110"), -- 0.4 + -0.6 = -0.2
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111011001100110011001101000"), -- -3 + 3.9 = 0.9
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000101001100110011001100110"), -- -3.3 + -1.9 = -5.2
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000110011001100110011001101"), -- 2.9 + 3.5 = 6.4
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111000110011001100110011010"), -- 0.6 + -0 = 0.6
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000010100110011001100110011"), -- -1.2 + -2.1 = -3.3
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111110110011001100110011010"), -- 0.5 + 1.2 = 1.7
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000010001100110011001100110"), -- -0.5 + 3.6 = 3.1
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000000001100110011001100110"), -- 2.6 + -0.5 = 2.1
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000101011001100110011001101"), -- -3.5 + -1.9 = -5.4
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000011110011001100110011010"), -- -2.9 + -1 = -3.9
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111110111111111111111111111111"), -- 0.4 + -0.9 = -0.5
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000110011001100110011010"), -- -3.8 + 1.4 = -2.4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000111100000000000000000000"), -- -3.8 + -3.7 = -7.5
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111000000000000000000000000"), -- -3 + 3.5 = 0.5
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000011011001100110011001100"), -- -2.8 + -0.9 = -3.7
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000010001100110011001100110"), -- 0.6 + 2.5 = 3.1
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000011100110011001100110011"), -- 3.7 + 0.1 = 3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000111010011001100110011010"), -- -3.9 + -3.4 = -7.3
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111110110011001100110011001110"), -- -0.7 + 1.1 = 0.4
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000100001100110011001100111"), -- -3.9 + -0.3 = -4.2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000000001100110011001100110"), -- 0.2 + 1.9 = 2.1
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"11000000000000000000000000000000"), -- -3.7 + 1.7 = -2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111101100110011001100110011"), -- -2.5 + 1.1 = -1.4
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0.6 + -0.3 = 0.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000001100110011001100110011"), -- -3.5 + 0.7 = -2.8
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111110110011001100110011010"), -- -2.2 + 3.9 = 1.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"10111111000000000000000000000000"), -- -3.6 + 3.1 = -0.5
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111110011001100110011001101"), -- -1.2 + -0.4 = -1.6
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111110110011001100110011001110"), -- -0.8 + 1.2 = 0.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000100101100110011001100110"), -- -1.1 + -3.6 = -4.7
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000011110011001100110011010"), -- 2.5 + 1.4 = 3.9
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000001011001100110011001101"), -- -0.7 + 3.4 = 2.7
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111001100110011001100110000"), -- 3.1 + -2.4 = 0.7
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000101000110011001100110011"), -- 1.6 + 3.5 = 5.1
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111110110011001100110011001100"), -- 1.5 + -1.1 = 0.4
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"00111111111001100110011001100111"), -- -1.9 + 3.7 = 1.8
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000001011001100110011001101"), -- -2.7 + -0 = -2.7
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00111111100110011001100110011010"), -- -1.3 + 2.5 = 1.2
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000110011001100110011001101"), -- -3 + -3.4 = -6.4
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"11000000000011001100110011001101"), -- -3 + 0.8 = -2.2
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000000011001100110011001100"), -- 2.6 + -0.4 = 2.2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000000001100110011001100110"), -- -1.1 + 3.2 = 2.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000100000000000000000000000"), -- -1.2 + -2.8 = -4
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110110011001100110011010"), -- 3.2 + 3.6 = 6.8
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111110110011001100110011010"), -- -2.1 + 3.8 = 1.7
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000101110011001100110011010"), -- -2 + -3.8 = -5.8
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000000001100110011001100110"), -- 0.9 + -3 = -2.1
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111010011001100110011001100"), -- -2 + 2.8 = 0.8
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000001100110011001100110011"), -- -0.5 + 3.3 = 2.8
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000001011001100110011001101"), -- -2.4 + -0.3 = -2.7
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000100000000000000000000000"), -- 1.6 + 2.4 = 4
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000100100000000000000000000"), -- -2.7 + -1.8 = -4.5
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"01000000000000000000000000000000"), -- 3.9 + -1.9 = 2
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001001100110011001100110"), -- 2.6 + -0 = 2.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000010100110011001100110011"), -- 1.5 + 1.8 = 3.3
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000010001100110011001100110"), -- 1.6 + 1.5 = 3.1
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000001000000000000000000000"), -- -1.5 + -1 = -2.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001000000000000000000000"), -- 2.5 + -0 = 2.5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000001100110011001100110011"), -- -0.7 + -2.1 = -2.8
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000000000000000000000000"), -- -3.4 + 1.4 = -2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000011011001100110011001100"), -- -1.1 + -2.6 = -3.7
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111100110011001100110011001"), -- -1.1 + 2.3 = 1.2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111110000000000000000000000"), -- 0.2 + 1.3 = 1.5
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111010011001100110011001100"), -- 1 + -1.8 = -0.8
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000101000000000000000000000"), -- -1.9 + -3.1 = -5
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111000000000000000000000000"), -- 3.2 + -2.7 = 0.5
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001100110011001100110011"), -- 3 + -0.2 = 2.8
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011110011001100110011001"), -- -0.1 + -3.8 = -3.9
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000011001100110011001101"), -- 0.2 + 2 = 2.2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000010100110011001100110011"), -- 0.7 + 2.6 = 3.3
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111100011001100110011001101"), -- -3 + 1.9 = -1.1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000001000000000000000000000"), -- 0.6 + 1.9 = 2.5
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000100001100110011001100110"), -- -1.4 + -2.8 = -4.2
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111011001100110011001100100"), -- 2.7 + -3.6 = -0.9
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111011001100110011001100110"), -- 1.5 + -0.6 = 0.9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000110100110011001100110100"), -- 2.9 + 3.7 = 6.6
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111001100110011001100110011"), -- -0.7 + -0 = -0.7
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111010011001100110011001110"), -- -2.7 + 1.9 = -0.8
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"00111101110011001100110011001110"), -- 0.3 + -0.2 = 0.1
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"00111111101100110011001100110100"), -- 2.9 + -1.5 = 1.4
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000000100110011001100110011"), -- 2 + 0.3 = 2.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001100110011001100110011"), -- -0.2 + -2.6 = -2.8
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"10111111111001100110011001100110"), -- 0.7 + -2.5 = -1.8
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000010011001100110011001101"), -- -2.7 + -0.5 = -3.2
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000110111001100110011001100"), -- -3.8 + -3.1 = -6.9
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111111010011001100110011001101"), -- -1 + 0.2 = -0.8
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000101111001100110011001101"), -- -3.5 + -2.4 = -5.9
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000010000000000000000000000"), -- -1.6 + -1.4 = -3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111101100110011001100110011"), -- -2.5 + 1.1 = -1.4
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000000011001100110011001101"), -- 2.5 + -0.3 = 2.2
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111110011001100110011001101"), -- 1.6 + -0 = 1.6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111110110011001100110011001100"), -- -1.4 + 1.8 = 0.4
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000100101100110011001100110"), -- -3.2 + -1.5 = -4.7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000000100110011001100110100"), -- 3.4 + -1.1 = 2.3
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111110000000000000000000000"), -- -2 + 3.5 = 1.5
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000010001100110011001100110"), -- -0.9 + -2.2 = -3.1
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111101001100110011001100110"), -- 1.4 + -0.1 = 1.3
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011000000000000000000000"), -- 0.3 + -3.8 = -3.5
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000111000000000000000000000"), -- -3.7 + -3.3 = -7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000010100110011001100110011"), -- 3.7 + -0.4 = 3.3
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000110001100110011001100110"), -- -2.7 + -3.5 = -6.2
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000011001100110011001100110"), -- 2.7 + 0.9 = 3.6
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111101100110011001100110011"), -- 0.5 + -1.9 = -1.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000101011001100110011001100"), -- -1.8 + -3.6 = -5.4
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111101100110011001100110011"), -- -1.3 + -0.1 = -1.4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000101010011001100110011010"), -- -3.8 + -1.5 = -5.3
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111111110110011001100110011001"), -- 1.4 + -3.1 = -1.7
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111101100110011001100110100"), -- 2.4 + -1 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111111110000000000000000000000"), -- 0.8 + -2.3 = -1.5
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111110100110011001100110011000"), -- 1.7 + -2 = -0.3
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000010001100110011001100110"), -- -0.9 + -2.2 = -3.1
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010011001100110011001101"), -- 0.2 + 3 = 3.2
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001100110011001100110011"), -- -0.1 + -2.7 = -2.8
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000101101100110011001100110"), -- -3 + -2.7 = -5.7
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00111111000000000000000000000000"), -- -2.6 + 3.1 = 0.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111110100110011001100110011000"), -- -3.2 + 3.5 = 0.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000000100110011001100110100"), -- 0.6 + -2.9 = -2.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000010100110011001100110011"), -- 2.1 + 1.2 = 3.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000111000110011001100110100"), -- 3.4 + 3.7 = 7.1
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111111001100110011001100110011"), -- -1 + 0.3 = -0.7
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000100000110011001100110011"), -- -3.4 + -0.7 = -4.1
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100000000000000000000000"), -- 0.1 + -1.1 = -1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001000000000000000000000"), -- 2.5 + -0 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000001000000000000000000000"), -- -0.9 + -1.6 = -2.5
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000100011001100110011001101"), -- 1.2 + 3.2 = 4.4
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000000110011001100110011010"), -- 2 + 0.4 = 2.4
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"10111111000110011001100110011100"), -- -2.9 + 2.3 = -0.6
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000010110011001100110011010"), -- 1.1 + 2.3 = 3.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"10111111110110011001100110011001"), -- -1.8 + 0.1 = -1.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000010001100110011001100110"), -- 1.1 + 2 = 3.1
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000110110011001100110011010"), -- -3.3 + -3.5 = -6.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000100101100110011001100110"), -- 3.7 + 1 = 4.7
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111110000000000000000000000"), -- -0.3 + 1.8 = 1.5
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111111100110011001100110100"), -- 0.8 + 1.1 = 1.9
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111110110011001100110011001100"), -- 1 + -1.4 = -0.4
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000100010011001100110011010"), -- -1.6 + -2.7 = -4.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111111110011001100110011001110"), -- 2.1 + -3.7 = -1.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"00111110100110011001100110011000"), -- 3.3 + -3 = 0.3
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111110100110011001100110011000"), -- 1.6 + -1.9 = -0.3
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000010110011001100110011010"), -- -1.4 + -2 = -3.4
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111001100110011001100110100"), -- -1 + 1.7 = 0.7
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000100001100110011001100110"), -- -2.6 + -1.6 = -4.2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000101101100110011001100110"), -- 2.4 + 3.3 = 5.7
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000101000110011001100110011"), -- -3.8 + -1.3 = -5.1
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111101001100110011001100110"), -- 0.3 + 1 = 1.3
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111111111100110011001100110100"), -- -2.7 + 0.8 = -1.9
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"10111110110011001100110011001100"), -- -1.8 + 1.4 = -0.4
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000100111001100110011001101"), -- 3.3 + 1.6 = 4.9
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000101000110011001100110100"), -- -2.2 + -2.9 = -5.1
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101110011001100110011010"), -- 2.8 + 3 = 5.8
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111000000000000000000000010"), -- -2.4 + 1.9 = -0.5
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000101100000000000000000000"), -- -2.3 + -3.2 = -5.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111111001100110011001100110010"), -- 1.9 + -1.2 = 0.7
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000100010011001100110011010"), -- -1.2 + -3.1 = -4.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000101100110011001100110011"), -- -3.5 + -2.1 = -5.6
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000100001100110011001100110"), -- -3.2 + -1 = -4.2
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111110111111111111111111111100"), -- -1.6 + 2.1 = 0.5
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111111111100110011001100110011"), -- -2.3 + 0.4 = -1.9
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111111001100110011001100110011"), -- 1.5 + -0.8 = 0.7
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111111110110011001100110011010"), -- 3.5 + -1.8 = 1.7
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111110100110011001100110011100"), -- 1.3 + -1.6 = -0.3
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111101001100110011001100111"), -- -2.4 + 1.1 = -1.3
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000101100000000000000000000"), -- -3 + -2.5 = -5.5
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000001011001100110011001101"), -- 1.1 + 1.6 = 2.7
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000100111001100110011001101"), -- -3 + -1.9 = -4.9
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"10111110100110011001100110011000"), -- 1.8 + -2.1 = -0.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111110110011001100110011001101"), -- -0.2 + -0.2 = -0.4
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111110000000000000000000000"), -- -2 + 3.5 = 1.5
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000001100110011001100110011"), -- -1.9 + -0.9 = -2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111000000000000000000000000"), -- 0 + 0.5 = 0.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000101000000000000000000000"), -- -3.2 + -1.8 = -5
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001100110011001100110011"), -- 3 + -0.2 = 2.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111110100110011001100110011000"), -- -2.8 + 2.5 = -0.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000011000000000000000000000"), -- -0.2 + -3.3 = -3.5
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111101001100110011001101000"), -- 3.4 + -2.1 = 1.3
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000000000100110011001100110100"), -- -2.9 + 0.6 = -2.3
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111111001100110011001100110"), -- 0.8 + 1 = 1.8
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000000000000000000000000000"), -- -0.7 + -1.3 = -2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111001100110011001100110011"), -- 0 + 0.7 = 0.7
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000011001100110011001100110"), -- -0.9 + -2.7 = -3.6
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000000000000000000000000000"), -- 1.6 + 0.4 = 2
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000010100110011001100110011"), -- -3.6 + 0.3 = -3.3
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"10111111110011001100110011001100"), -- 0.5 + -2.1 = -1.6
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111000000000000000000000000"), -- 1.6 + -1.1 = 0.5
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111100110011001100110011010"), -- 3.3 + -2.1 = 1.2
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000101111001100110011001101"), -- -3.4 + -2.5 = -5.9
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000000000000000000000000000"), -- 1.9 + 0.1 = 2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000000000000000000000000000"), -- -0.3 + -1.7 = -2
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"10111111000110011001100110011000"), -- 1.5 + -2.1 = -0.6
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000011000000000000000000000"), -- 3.4 + 0.1 = 3.5
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"10111111011001100110011001101000"), -- -2.2 + 1.3 = -0.9
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000011110011001100110011001"), -- 1.3 + 2.6 = 3.9
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000100000000000000000000000"), -- 0.6 + 3.4 = 4
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111110110011001100110011010"), -- -0.5 + 2.2 = 1.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111101110011001100110011010000"), -- 1.1 + -1 = 0.1
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111101110011001100110011010000"), -- 0.8 + -0.7 = 0.1
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"10111110100110011001100110100000"), -- -2.4 + 2.1 = -0.3
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"10111111101100110011001100110011"), -- -1.9 + 0.5 = -1.4
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111100011001100110011001101"), -- -2.7 + 1.6 = -1.1
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000111010011001100110011010"), -- 3.4 + 3.9 = 7.3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101100110011001100110011"), -- 2.6 + 3 = 5.6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000000110011001100110011010"), -- 0.8 + -3.2 = -2.4
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000011110011001100110011010"), -- 1.5 + 2.4 = 3.9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000101010011001100110011010"), -- 2.9 + 2.4 = 5.3
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000111010011001100110011010"), -- -3.9 + -3.4 = -7.3
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000100001100110011001100111"), -- 3.9 + 0.3 = 4.2
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000001100110011001100110011"), -- 0.9 + 1.9 = 2.8
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001011001100110011001101"), -- 2.7 + -0 = 2.7
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000000100110011001100110011"), -- 2.5 + -0.2 = 2.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000010110011001100110011010"), -- -1.2 + -2.2 = -3.4
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111110100110011001100110011000"), -- 3.4 + -3.7 = -0.3
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000101110011001100110011010"), -- 2.5 + 3.3 = 5.8
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000110101100110011001100110"), -- -2.9 + -3.8 = -6.7
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000100001100110011001100111"), -- -0.3 + -3.9 = -4.2
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111111110110011001100110011001"), -- -2.1 + 0.4 = -1.7
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000111001100110011001100110"), -- -3.3 + -3.9 = -7.2
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111110000000000000000000000"), -- 1.5 + -0 = 1.5
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111110011001100110011001100"), -- -0.3 + -1.3 = -1.6
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111110010011001100110011010000"), -- -2.7 + 2.5 = -0.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111110110011001100110011001100"), -- -0.7 + 0.3 = -0.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000011100110011001100110011"), -- -1.8 + -2 = -3.8
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"10111110100110011001100110100000"), -- -3.9 + 3.6 = -0.3
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000011100110011001100110100"), -- 1.1 + 2.7 = 3.8
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000001001100110011001100110"), -- 0.5 + -3.1 = -2.6
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000101011001100110011001101"), -- 3.4 + 2 = 5.4
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000100110011001100110011010"), -- 2.4 + 2.4 = 4.8
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000000100110011001100110011"), -- 1.5 + -3.8 = -2.3
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111110011001100110011001101"), -- -0.8 + -0.8 = -1.6
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111110010011001100110011010000"), -- -3 + 2.8 = -0.2
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111000000000000000000000000"), -- -3.4 + 3.9 = 0.5
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000000011001100110011001101"), -- -1.8 + -0.4 = -2.2
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111110100110011001100110011000"), -- -3.3 + 3.6 = 0.3
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000101111001100110011001101"), -- -2.4 + -3.5 = -5.9
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000000001100110011001100110"), -- -0.5 + -1.6 = -2.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111110100110011001100110011010"), -- 0 + -0.3 = -0.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000101000110011001100110011"), -- -3.6 + -1.5 = -5.1
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010001100110011001100111"), -- -0.3 + 3.4 = 3.1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111111101001100110011001100110"), -- 2.1 + -0.8 = 1.3
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000001110011001100110011010"), -- 1.3 + 1.6 = 2.9
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111111001100110011001100111"), -- -2.4 + 0.6 = -1.8
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000000011001100110011001100"), -- 1.1 + -3.3 = -2.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011000000000000000000000"), -- -0.2 + 3.7 = 3.5
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000110100000000000000000000"), -- 3.6 + 2.9 = 6.5
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000010011001100110011001101"), -- -2.5 + -0.7 = -3.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111110110011001100110011001"), -- 2.8 + -1.1 = 1.7
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"), -- -3.1 + 3.1 = 0
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"00111111011001100110011001101000"), -- 3.7 + -2.8 = 0.9
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000100110011001100110011010"), -- -1.6 + -3.2 = -4.8
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000101010011001100110011010"), -- -2.6 + -2.7 = -5.3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111111100110011001100110011"), -- -2.5 + 0.6 = -1.9
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000000001001100110011001100111"), -- -2.7 + 0.1 = -2.6
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111110010011001100110011000000"), -- 2.9 + -3.1 = -0.2
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001011001100110011001101"), -- 2.9 + -0.2 = 2.7
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000010100110011001100110011"), -- -0.7 + -2.6 = -3.3
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100001100110011001100110"), -- 1.1 + 3.1 = 4.2
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111110100110011001100110011000"), -- -3.3 + 3.6 = 0.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111110010011001100110011001100"), -- -0.6 + 0.8 = 0.2
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000100001100110011001100110"), -- -1.8 + -2.4 = -4.2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"00111110100110011001100110011000"), -- 2 + -1.7 = 0.3
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111000110011001100110011000"), -- 3 + -2.4 = 0.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110010011001100110011010"), -- 2.7 + 3.6 = 6.3
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000000001100110011001100111"), -- -0.4 + -1.7 = -2.1
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000000000000000000000000000"), -- -0.1 + -1.9 = -2
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000001000000000000000000000"), -- -1 + -1.5 = -2.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000001110011001100110011010"), -- -3.2 + 0.3 = -2.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000010011001100110011001101"), -- 3 + 0.2 = 3.2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111110110011001100110011001100"), -- -0.3 + 0.7 = 0.4
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100100110011001100110011"), -- 1.5 + 3.1 = 4.6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000100010011001100110011010"), -- -1.4 + -2.9 = -4.3
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100110011001100110011010"), -- -0.1 + -1.1 = -1.2
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000001001100110011001100110"), -- 0.5 + -3.1 = -2.6
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000100010011001100110011010"), -- -2.6 + -1.7 = -4.3
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"10111110100110011001100110011000"), -- -2.7 + 2.4 = -0.3
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000000000000000000000000000"), -- 0.3 + 1.7 = 2
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000011110011001100110011010"), -- -2.7 + -1.2 = -3.9
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000101010011001100110011010"), -- -1.7 + -3.6 = -5.3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"10111111110011001100110011001101"), -- 0.9 + -2.5 = -1.6
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111101100110011001100110011"), -- -0.5 + -0.9 = -1.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000110011001100110011001101"), -- -3.7 + -2.7 = -6.4
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000000000000000000000000000"), -- -1.7 + 3.7 = 2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111100000000000000000000000"), -- -2.5 + 1.5 = -1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000011001100110011001100110"), -- 2.1 + 1.5 = 3.6
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"10111111010011001100110011001100"), -- 2.4 + -3.2 = -0.8
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000011000000000000000000000"), -- -0.1 + 3.6 = 3.5
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000001100110011001100110011"), -- 2.6 + 0.2 = 2.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000101110011001100110011010"), -- 3.8 + 2 = 5.8
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000100001100110011001100110"), -- -0.5 + -3.7 = -4.2
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111100000000000000000000000"), -- -1.3 + 2.3 = 1
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111110010011001100110011001100"), -- 1 + -0.8 = 0.2
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"10111101110011001100110011000000"), -- -2.8 + 2.7 = -0.0999999
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111110000000000000000000000"), -- 0 + -1.5 = -1.5
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"10111110100110011001100110011000"), -- -3.3 + 3 = -0.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000100000110011001100110011"), -- 3.4 + 0.7 = 4.1
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000001001100110011001100110"), -- 3.6 + -1 = 2.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"), -- -2 + 2 = 0
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111110010011001100110011010000"), -- 1.2 + -1 = 0.2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011011001100110011001101"), -- 0.2 + 3.5 = 3.7
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000101011001100110011001101"), -- 2.7 + 2.7 = 5.4
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000001001100110011001100110"), -- -1.6 + -1 = -2.6
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111001100110011001100110011"), -- -0.2 + 0.9 = 0.7
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000001000000000000000000000"), -- 0.9 + 1.6 = 2.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111111110110011001100110011010"), -- 2.5 + -0.8 = 1.7
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101011001100110011001101"), -- 3.2 + 2.2 = 5.4
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111111110000000000000000000001"), -- -2.4 + 0.9 = -1.5
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111101100110011001100110100"), -- -2.5 + 3.9 = 1.4
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100011001100110011001101"), -- 0.9 + 3.5 = 4.4
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000000000000000000000000000"), -- -1.4 + -0.6 = -2
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000111010011001100110011010"), -- -3.5 + -3.8 = -7.3
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111110110011001100110011010"), -- -1.4 + -0.3 = -1.7
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111010011001100110011010000"), -- 2.1 + -2.9 = -0.8
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111100110011001100110011001"), -- 0.2 + -1.4 = -1.2
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111110110011001100110011001100"), -- 0.9 + -0.5 = 0.4
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111110011001100110011001100"), -- -0.7 + 2.3 = 1.6
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111110010011001100110011010000"), -- 2.1 + -2.3 = -0.2
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000011011001100110011001101"), -- -3.2 + -0.5 = -3.7
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101011001100110011001101"), -- 2.9 + 2.5 = 5.4
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000100100110011001100110011"), -- 3.8 + 0.8 = 4.6
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101011001100110011001101"), -- -3.8 + -1.6 = -5.4
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000111010011001100110011010"), -- 3.4 + 3.9 = 7.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000011001100110011001100111"), -- -1.2 + -2.4 = -3.6
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000010100110011001100110011"), -- 1.2 + 2.1 = 3.3
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000100110011001100110100"), -- -0.1 + 2.4 = 2.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000111000000000000000000000"), -- -3.6 + -3.4 = -7
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000110000110011001100110011"), -- 2.8 + 3.3 = 6.1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000100001100110011001100110"), -- 2.1 + 2.1 = 4.2
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111100110011001100110011010"), -- -0.8 + -0.4 = -1.2
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000110011001100110011001101"), -- 3 + 3.4 = 6.4
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111101110011001100110011000000"), -- 2.1 + -2 = 0.0999999
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000000001100110011001100111"), -- -1.7 + -0.4 = -2.1
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111101100110011001100110010"), -- 1.2 + -2.6 = -1.4
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111100011001100110011001100"), -- -1.7 + 2.8 = 1.1
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010001100110011001100111"), -- -0.3 + 3.4 = 3.1
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000011001100110011001100110"), -- -1.6 + -2 = -3.6
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100000000000000000000000"), -- 0.1 + -1.1 = -1
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000001000000000000000000000"), -- -2.5 + -0 = -2.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000011011001100110011001101"), -- -3.2 + -0.5 = -3.7
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000011100110011001100110011"), -- -3 + -0.8 = -3.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000011100110011001100110011"), -- 0 + -3.8 = -3.8
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111110010011001100110011010000"), -- 2.7 + -2.5 = 0.2
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100100000000000000000000"), -- 1.4 + 3.1 = 4.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000101111001100110011001101"), -- -3.2 + -2.7 = -5.9
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111110011001100110011001101"), -- -1.6 + -0 = -1.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111110010011001100110011010000"), -- 2.7 + -2.9 = -0.2
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000000011001100110011001101"), -- 1.1 + 1.1 = 2.2
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111111100011001100110011001101"), -- 0.9 + -2 = -1.1
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000100011001100110011001101"), -- 3.4 + 1 = 4.4
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000100111001100110011001101"), -- 3.2 + 1.7 = 4.9
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000001011001100110011001100"), -- -0.1 + -2.6 = -2.7
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000000001100110011001100110"), -- 1.5 + 0.6 = 2.1
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111110011001100110011001110"), -- 3.7 + -2.1 = 1.6
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000000001110011001100110011010"), -- 3.7 + -0.8 = 2.9
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000001100110011001100110100"), -- -2.4 + -0.4 = -2.8
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000101100000000000000000000"), -- 2.1 + 3.4 = 5.5
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111110110011001100110011010"), -- -0.5 + -1.2 = -1.7
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000110001100110011001100110"), -- -3.7 + -2.5 = -6.2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000101100000000000000000000"), -- -2.5 + -3 = -5.5
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000010100110011001100110011"), -- 0.2 + -3.5 = -3.3
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"), -- 0.4 + -0.4 = 0
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111101001100110011001100111"), -- -0.9 + 2.2 = 1.3
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111110010011001100110011001000"), -- 1.7 + -1.9 = -0.2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000000110011001100110011010"), -- -1.1 + 3.5 = 2.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111111011001100110011001101000"), -- -3.7 + 2.8 = -0.9
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000110100110011001100110100"), -- 2.7 + 3.9 = 6.6
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"10111111101100110011001100110100"), -- -3.7 + 2.3 = -1.4
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000010100110011001100110011"), -- 3.8 + -0.5 = 3.3
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001110011001100110011010"), -- 2.9 + -0 = 2.9
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000100111001100110011001100"), -- -3.6 + -1.3 = -4.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"10111110110011001100110011010000"), -- 2.8 + -3.2 = -0.4
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111111100110011001100110010"), -- -0.7 + 2.6 = 1.9
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000100001100110011001100110"), -- 3.5 + 0.7 = 4.2
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111111000110011001100110011000"), -- -1.5 + 2.1 = 0.6
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111101110011001100110011000000"), -- -2.5 + 2.6 = 0.0999999
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111110000000000000000000001"), -- -3.4 + 1.9 = -1.5
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000110100110011001100110011"), -- -3.8 + -2.8 = -6.6
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101000110011001100110100"), -- 2.9 + 2.2 = 5.1
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000100000000000000000000000"), -- -2.6 + -1.4 = -4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000000100110011001100110011"), -- -3.3 + 1 = -2.3
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111111100011001100110011001100"), -- -1.8 + 0.7 = -1.1
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111110100110011001100110011000"), -- -2.1 + 1.8 = -0.3
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"00111111011001100110011001100111"), -- 1.1 + -0.2 = 0.9
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000001001100110011001100111"), -- 0.4 + 2.2 = 2.6
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111110010011001100110011000000"), -- 2.9 + -3.1 = -0.2
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000100001100110011001100110"), -- -1.7 + -2.5 = -4.2
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000010100110011001100110100"), -- 3.9 + -0.6 = 3.3
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000001011001100110011001101"), -- -0.3 + -2.4 = -2.7
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000000011001100110011001101"), -- 1.8 + 0.4 = 2.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000010100110011001100110011"), -- -0.5 + 3.8 = 3.3
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000110000110011001100110100"), -- -3.9 + -2.2 = -6.1
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"00111110110011001100110011010000"), -- -2.6 + 3 = 0.4
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100110011001100110011010"), -- -0.1 + -1.1 = -1.2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000001000000000000000000000"), -- -1.1 + -1.4 = -2.5
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000101100000000000000000000"), -- 1.6 + 3.9 = 5.5
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000010100110011001100110011"), -- -3.3 + -0 = -3.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000100000110011001100110011"), -- 3.4 + 0.7 = 4.1
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000001110011001100110011010"), -- 3.4 + -0.5 = 2.9
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"), -- -1.4 + 1.4 = 0
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000110100000000000000000000"), -- -2.6 + -3.9 = -6.5
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000010000000000000000000000"), -- 0.3 + -3.3 = -3
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000011100110011001100110100"), -- 2.7 + 1.1 = 3.8
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111111011001100110011001101000"), -- -2 + 2.9 = 0.9
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111001100110011001100110100"), -- 0.4 + -1.1 = -0.7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000101110011001100110011010"), -- 3.4 + 2.4 = 5.8
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000101110011001100110011010"), -- -3.3 + -2.5 = -5.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000000000011001100110011001100"), -- -2.8 + 0.6 = -2.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000001000000000000000000000"), -- -0.9 + -1.6 = -2.5
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000000000000000000000000000"), -- 1.6 + 0.4 = 2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111101110011001100110011000000"), -- -1.2 + 1.3 = 0.0999999
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111111000000000000000000000000"), -- 2.2 + -2.7 = -0.5
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111111101100110011001100110011"), -- -1.6 + 0.2 = -1.4
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111100000000000000000000000"), -- 3.5 + -2.5 = 1
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111110011001100110011001110"), -- 1.8 + -3.4 = -1.6
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111000110011001100110011010"), -- 1.7 + -1.1 = 0.6
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000000110011001100110011010"), -- -0.4 + -2 = -2.4
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111110100110011001100110011000"), -- -3.2 + 3.5 = 0.3
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111100110011001100110011010"), -- -2.6 + 3.8 = 1.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000000001100110011001100110"), -- -0.9 + 3 = 2.1
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000000001100110011001100110"), -- -2.1 + -0 = -2.1
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000001001100110011001100110"), -- 1.5 + 1.1 = 2.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111101100110011001100110011"), -- -0.1 + 1.5 = 1.4
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000110001100110011001100110"), -- -2.4 + -3.8 = -6.2
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000101110011001100110011010"), -- -3.3 + -2.5 = -5.8
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000001100110011001100110011"), -- 2 + 0.8 = 2.8
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000011011001100110011001101"), -- 1.3 + 2.4 = 3.7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000101100000000000000000000"), -- 3.4 + 2.1 = 5.5
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"00111111000000000000000000000000"), -- 2.8 + -2.3 = 0.5
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011100110011001100110011"), -- 0.5 + 3.3 = 3.8
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000100111001100110011001101"), -- -1.4 + -3.5 = -4.9
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000001000000000000000000000"), -- -1.2 + -1.3 = -2.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000100000000000000000000000"), -- 0.4 + 3.6 = 4
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111111100110011001100110011010"), -- 1.7 + -0.5 = 1.2
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000011110011001100110011010"), -- -1.4 + -2.5 = -3.9
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000100101100110011001100110"), -- 3.2 + 1.5 = 4.7
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111110000000000000000000000"), -- -1.1 + -0.4 = -1.5
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000001100110011001100110011"), -- 3.3 + -0.5 = 2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000010000000000000000000000"), -- 0 + -3 = -3
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111111001100110011001100110"), -- 0.8 + 1 = 1.8
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110010011001100110011001101"), -- 0.2 + -0.4 = -0.2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111000110011001100110011010"), -- -0.3 + -0.3 = -0.6
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000101001100110011001100110"), -- 3.2 + 2 = 5.2
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100110011001100110011010"), -- 1.3 + 3.5 = 4.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111110110011001100110011010"), -- -0.3 + -1.4 = -1.7
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000101011001100110011001100"), -- 2.8 + 2.6 = 5.4
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111111100011001100110011001100"), -- -3.6 + 2.5 = -1.1
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000011011001100110011001100"), -- -0.9 + -2.8 = -3.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000111000110011001100110011"), -- -3.6 + -3.5 = -7.1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000001000000000000000000000"), -- -0.8 + 3.3 = 2.5
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000000011001100110011001101"), -- 0.7 + -2.9 = -2.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000010100110011001100110011"), -- -0.5 + -2.8 = -3.3
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111100110011001100110011010"), -- 3.9 + -2.7 = 1.2
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111001100110011001100110100"), -- -3.2 + 3.9 = 0.7
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000100010011001100110011010"), -- 3.5 + 0.8 = 4.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000000001001100110011001100110"), -- 2.1 + 0.5 = 2.6
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111111111100110011001100110100"), -- -3.7 + 1.8 = -1.9
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111100011001100110011001100"), -- -1.7 + 2.8 = 1.1
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111011001100110011001100100"), -- -2.4 + 3.3 = 0.9
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111010011001100110011001110"), -- -0.4 + 1.2 = 0.8
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000100111001100110011001100"), -- 1.3 + 3.6 = 4.9
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111111101001100110011001100110"), -- -3.1 + 1.8 = -1.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000011100110011001100110011"), -- 2.8 + 1 = 3.8
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111111100110011001100110010"), -- 1.7 + -3.6 = -1.9
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111101111111111111111111111"), -- -3.1 + 1.6 = -1.5
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111010011001100110011001100"), -- -2 + 1.2 = -0.8
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111101001100110011001100110"), -- -0.8 + -0.5 = -1.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000101110011001100110011010"), -- -3.6 + -2.2 = -5.8
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000010000000000000000000000"), -- -2.6 + -0.4 = -3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111101100110011001100110011"), -- -0.5 + -0.9 = -1.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000101000110011001100110011"), -- -1.8 + -3.3 = -5.1
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010011001100110011001101"), -- 0.2 + 3 = 3.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000100100000000000000000000"), -- -0.7 + -3.8 = -4.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000101000000000000000000000"), -- 1.9 + 3.1 = 5
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00111110100110011001100110011000"), -- -2.8 + 3.1 = 0.3
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000100100110011001100110011"), -- -1.1 + -3.5 = -4.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000100001100110011001100110"), -- 2.7 + 1.5 = 4.2
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111111101001100110011001100110"), -- 3.3 + -2 = 1.3
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001100110011001100110011"), -- 0.1 + 2.7 = 2.8
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111100110011001100110011010"), -- -3.2 + 2 = -1.2
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000000011001100110011001101"), -- 1.7 + -3.9 = -2.2
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101001100110011001100110"), -- -2.6 + -2.6 = -5.2
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111111111100110011001100110011"), -- 0.1 + -2 = -1.9
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000111000110011001100110100"), -- 3.9 + 3.2 = 7.1
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000000100110011001100110011"), -- 0.5 + 1.8 = 2.3
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000110010011001100110011010"), -- -3.3 + -3 = -6.3
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111111100110011001100110100"), -- -0.8 + -1.1 = -1.9
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011001100110011001100110"), -- 0.3 + 3.3 = 3.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000101011001100110011001101"), -- 2 + 3.4 = 5.4
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"), -- -3.5 + 3.5 = 0
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111110110011001100110011010000"), -- -2.3 + 2.7 = 0.4
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111111100110011001100110011010"), -- 3.2 + -2 = 1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111101110011001100110011001101"), -- 0 + 0.1 = 0.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000100110011001100110011010"), -- -1.2 + -3.6 = -4.8
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000011110011001100110011010"), -- 2 + 1.9 = 3.9
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"10111111100110011001100110011010"), -- 1.8 + -3 = -1.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111101001100110011001100111"), -- -0.2 + -1.1 = -1.3
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000010011001100110011001101"), -- -3.7 + 0.5 = -3.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000010100110011001100110011"), -- 3.2 + 0.1 = 3.3
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000010110011001100110011010"), -- -3.4 + -0 = -3.4
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111101001100110011001100110"), -- -0.5 + 1.8 = 1.3
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000000000001100110011001100111"), -- -2.2 + 0.1 = -2.1
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"), -- -1.9 + 1.9 = 0
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111111010011001100110011001101"), -- -1.5 + 0.7 = -0.8
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"00111111100000000000000000000000"), -- -2 + 3 = 1
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"), -- -1.5 + 1.5 = 0
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110001100110011001100110"), -- -3.3 + -2.9 = -6.2
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111110111111111111111111111110"), -- 0.8 + -1.3 = -0.5
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000110000000000000000000000"), -- 3.3 + 2.7 = 6
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"10111110110011001100110011010000"), -- -2.7 + 2.3 = -0.4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111110011001100110011001101"), -- 2.7 + -1.1 = 1.6
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000111100110011001100110100"), -- -3.9 + -3.7 = -7.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111011001100110011001100100"), -- 2.7 + -3.6 = -0.9
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111101110011001100110011100000"), -- 2.6 + -2.7 = -0.1
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111110000000000000000000000"), -- -1.3 + 2.8 = 1.5
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"00111111000000000000000000000000"), -- 3.7 + -3.2 = 0.5
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000110101100110011001100110"), -- 3.2 + 3.5 = 6.7
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000001011001100110011001101"), -- -0.8 + -1.9 = -2.7
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000101110011001100110011010"), -- -3 + -2.8 = -5.8
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111010011001100110011001101"), -- 0.1 + 0.7 = 0.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000110011001100110011001100"), -- -2.8 + -3.6 = -6.4
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111101001100110011001100110"), -- -0.5 + 1.8 = 1.3
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111010011001100110011001100"), -- 2 + -2.8 = -0.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111101001100110011001100110"), -- 1.4 + -0.1 = 1.3
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000101000110011001100110011"), -- 1.3 + 3.8 = 5.1
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"00111111101001100110011001100110"), -- 2.8 + -1.5 = 1.3
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111111001100110011001100110"), -- 1.4 + 0.4 = 1.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"00111111011001100110011001100100"), -- 3.8 + -2.9 = 0.9
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"00111101110011001100110011010000"), -- -1.9 + 2 = 0.1
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000100010011001100110011010"), -- 1.4 + 2.9 = 4.3
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000000000000000000000000000"), -- 3.5 + -1.5 = 2
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000101100110011001100110100"), -- -3.9 + -1.7 = -5.6
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111000110011001100110011010"), -- -1 + 1.6 = 0.6
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001110011001100110011010"), -- 2.9 + -0 = 2.9
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111101110011001100110011000000"), -- 2.2 + -2.3 = -0.0999999
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000011001100110011001100111"), -- 3.4 + 0.2 = 3.6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111111001100110011001100110"), -- -1.4 + -0.4 = -1.8
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000100100000000000000000000"), -- 1.7 + 2.8 = 4.5
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000110000000000000000000000"), -- -2.6 + -3.4 = -6
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111100000000000000000000000"), -- 1.6 + -0.6 = 1
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000101000000000000000000000"), -- 1.9 + 3.1 = 5
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111111101001100110011001100111"), -- -1.1 + 2.4 = 1.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111000000000000000000000000"), -- 0.6 + -0.1 = 0.5
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111110110011001100110011001100"), -- 1.4 + -1 = 0.4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111010011001100110011001110"), -- 2.7 + -1.9 = 0.8
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000000100110011001100110011"), -- 0.7 + 1.6 = 2.3
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000000000000000000000000000"), -- -0.7 + -1.3 = -2
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000110100110011001100110100"), -- -2.9 + -3.7 = -6.6
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111111100110011001100110011"), -- -2.5 + 0.6 = -1.9
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000101011001100110011001100"), -- 2.6 + 2.8 = 5.4
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111111001100110011001100110100"), -- -1.7 + 2.4 = 0.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000011011001100110011001100"), -- 1.1 + 2.6 = 3.7
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111100011001100110011001101"), -- -2.2 + 1.1 = -1.1
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000100000110011001100110011"), -- 2 + 2.1 = 4.1
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000010100110011001100110100"), -- 0.4 + 2.9 = 3.3
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000100100000000000000000000"), -- 1.9 + 2.6 = 4.5
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111011001100110011001101000"), -- -1.3 + 2.2 = 0.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101000000000000000000000"), -- 2.8 + 2.2 = 5
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000000001110011001100110011010"), -- 3.8 + -0.9 = 2.9
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000000000000000000000000000"), -- -1.9 + 3.9 = 2
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000001000000000000000000000"), -- 1.6 + 0.9 = 2.5
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000100111001100110011001101"), -- -2.7 + -2.2 = -4.9
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011110011001100110011010"), -- 0.6 + 3.3 = 3.9
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111101110011001100110011000000"), -- 3.2 + -3.3 = -0.0999999
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111110100110011001100110011000"), -- -1.4 + 1.1 = -0.3
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000010001100110011001100111"), -- -0.8 + 3.9 = 3.1
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111110110011001100110011010"), -- -0.3 + -1.4 = -1.7
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111111001100110011001100110011"), -- -1 + 0.3 = -0.7
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"10111111111001100110011001100110"), -- -1.9 + 0.1 = -1.8
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111010011001100110011001100"), -- -2 + 2.8 = 0.8
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000100010011001100110011010"), -- -2.7 + -1.6 = -4.3
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"), -- -3.7 + 3.7 = 0
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111101110011001100110011010000"), -- -0.9 + 1 = 0.1
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111100000000000000000000000"), -- -2.5 + 1.5 = -1
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000010011001100110011001100"), -- 1.8 + 1.4 = 3.2
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000000100110011001100110011"), -- 0.8 + -3.1 = -2.3
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001000000000000000000000"), -- 0.3 + -2.8 = -2.5
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000100100110011001100110100"), -- -3.4 + -1.2 = -4.6
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000011001100110011001100110"), -- -2.2 + -1.4 = -3.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000000011001100110011001101"), -- -1.3 + 3.5 = 2.2
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000101110011001100110011010"), -- 2.3 + 3.5 = 5.8
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111010011001100110011001100"), -- 1 + -1.8 = -0.8
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000101101100110011001100110"), -- 1.8 + 3.9 = 5.7
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000100000110011001100110011"), -- -0.4 + -3.7 = -4.1
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111101001100110011001100110"), -- 2.3 + -3.6 = -1.3
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111010011001100110011001100"), -- -2.8 + 2 = -0.8
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000010100110011001100110100"), -- 2.2 + 1.1 = 3.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000000011001100110011001100"), -- 0.6 + -2.8 = -2.2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000000110011001100110011001"), -- 0.7 + -3.1 = -2.4
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000001000000000000000000000"), -- 2.3 + 0.2 = 2.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000110011001100110011001101"), -- 3.5 + 2.9 = 6.4
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000101110011001100110011010"), -- -2 + -3.8 = -5.8
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111111100110011001100110100"), -- -0.2 + -1.7 = -1.9
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"10111111000110011001100110011000"), -- -3.3 + 2.7 = -0.6
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111101001100110011001100111"), -- 0.2 + 1.1 = 1.3
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"00111111101100110011001100110100"), -- 3.7 + -2.3 = 1.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111110110011001100110011001"), -- -3.3 + 1.6 = -1.7
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111111100011001100110011001110"), -- -2.9 + 1.8 = -1.1
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000100011001100110011001100"), -- -3.1 + -1.3 = -4.4
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000011110011001100110011010"), -- 2.2 + 1.7 = 3.9
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111110110011001100110011010"), -- -2.9 + 1.2 = -1.7
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"10111111100110011001100110011010"), -- 1 + -2.2 = -1.2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111101100110011001100110100"), -- -1.1 + -0.3 = -1.4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000011110011001100110011010"), -- 2.7 + 1.2 = 3.9
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000011001100110011001100110"), -- 1.7 + 1.9 = 3.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110111001100110011001100"), -- 3.3 + 3.6 = 6.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111001100110011001100110100"), -- -0.3 + -0.4 = -0.7
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"00111110110011001100110011010000"), -- 3.2 + -2.8 = 0.4
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000000100110011001100110011"), -- 3.3 + -1 = 2.3
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111110100110011001100110011000"), -- -1.9 + 1.6 = -0.3
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000101000110011001100110100"), -- -3.9 + -1.2 = -5.1
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111101110011001100110011001110"), -- -0.3 + 0.2 = -0.1
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000010100110011001100110100"), -- -0.4 + -2.9 = -3.3
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111110110011001100110011001000"), -- -3.4 + 3.8 = 0.4
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000010001100110011001100110"), -- -0.3 + -2.8 = -3.1
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000001110011001100110011010"), -- -2 + -0.9 = -2.9
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111110000000000000000000000"), -- -2.7 + 1.2 = -1.5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000010001100110011001100110"), -- -0.7 + 3.8 = 3.1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000011011001100110011001101"), -- -0.7 + -3 = -3.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000011110011001100110011001"), -- -3.6 + -0.3 = -3.9
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111110110011001100110011001100"), -- 0.9 + -1.3 = -0.4
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111111001100110011001100111"), -- -2.4 + 0.6 = -1.8
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000100001100110011001100110"), -- -3.5 + -0.7 = -4.2
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111101100110011001100110010"), -- -2.4 + 3.8 = 1.4
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111100000000000000000000000"), -- 0.8 + 0.2 = 1
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011011001100110011001101"), -- -0.2 + -3.5 = -3.7
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000100000000000000000000000"), -- -1.4 + -2.6 = -4
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000000100110011001100110011"), -- 3.8 + -1.5 = 2.3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111111000110011001100110011001"), -- 0.9 + -0.3 = 0.6
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111111000110011001100110011100"), -- -1.8 + 2.4 = 0.6
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"10111111010011001100110011001100"), -- -3.2 + 2.4 = -0.8
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000001000000000000000000000"), -- -0.9 + -1.6 = -2.5
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111110111111111111111111111110"), -- -0.8 + 1.3 = 0.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000110000110011001100110011"), -- 3.5 + 2.6 = 6.1
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111111100110011001100110100"), -- 0.7 + 1.2 = 1.9
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"10111110010011001100110011010000"), -- -2.3 + 2.1 = -0.2
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000110101100110011001100110"), -- 2.9 + 3.8 = 6.7
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000111000110011001100110011"), -- -3.5 + -3.6 = -7.1
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"11000000001001100110011001100111"), -- -3.4 + 0.8 = -2.6
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111000110011001100110011010"), -- 2.5 + -1.9 = 0.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000000011001100110011001101"), -- 1.5 + -3.7 = -2.2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000011001100110011001100111"), -- -1.2 + -2.4 = -3.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111111100110011001100110011"), -- 2 + -0.1 = 1.9
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111011001100110011001101000"), -- -3 + 3.9 = 0.9
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"00111111000000000000000000000000"), -- 3.3 + -2.8 = 0.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"00111111001100110011001100110100"), -- 3.5 + -2.8 = 0.7
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000110101100110011001100110"), -- 3.3 + 3.4 = 6.7
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000000001100110011001100111"), -- 0.8 + -2.9 = -2.1
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111111111111111111111111111"), -- 1.6 + -3.6 = -2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000001100110011001100110011"), -- 3.2 + -0.4 = 2.8
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000000000000000000000000000"), -- -3.2 + 1.2 = -2
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000010000000000000000000000"), -- 0.4 + 2.6 = 3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111011001100110011001100111"), -- 0.7 + -1.6 = -0.9
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000000100110011001100110011"), -- -0.4 + -1.9 = -2.3
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"10111111100011001100110011001100"), -- -3.8 + 2.7 = -1.1
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111111100110011001100110100"), -- 1.7 + 0.2 = 1.9
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000101110011001100110011010"), -- 3.5 + 2.3 = 5.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000011110011001100110011010"), -- 1.4 + 2.5 = 3.9
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111000000000000000000000000"), -- 2.6 + -2.1 = 0.5
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111111001100110011001100110"), -- -0.8 + 2.6 = 1.8
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"10111111111100110011001100110011"), -- 0.6 + -2.5 = -1.9
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000101101100110011001100110"), -- 2 + 3.7 = 5.7
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111001100110011001100110010"), -- 0.6 + -1.3 = -0.7
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000000001100110011001100110"), -- 2.1 + -0 = 2.1
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111101110011001100110011000000"), -- -2 + 2.1 = 0.0999999
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111101001100110011001100110"), -- 2.3 + -1 = 1.3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111110010011001100110011001100"), -- 0.7 + -0.5 = 0.2
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000000001100110011001100110"), -- -0.4 + 2.5 = 2.1
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000011100110011001100110011"), -- 3.8 + -0 = 3.8
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111000110011001100110011000"), -- 2.2 + -2.8 = -0.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000110011001100110011001100"), -- 3.3 + 3.1 = 6.4
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"10111101110011001100110011010000"), -- -1.4 + 1.3 = -0.1
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000100010011001100110011010"), -- -2.9 + -1.4 = -4.3
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000111011001100110011001101"), -- 3.5 + 3.9 = 7.4
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111001100110011001100110100"), -- 3.2 + -2.5 = 0.7
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000000100110011001100110011"), -- -1.3 + 3.6 = 2.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101000110011001100110011"), -- 2.1 + 3 = 5.1
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000000110011001100110011010"), -- 1.4 + -3.8 = -2.4
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111110110011001100110011001110"), -- -1.2 + 0.8 = -0.4
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000001001100110011001100111"), -- 2.2 + 0.4 = 2.6
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111111001100110011001100110"), -- -0.4 + -1.4 = -1.8
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000101110011001100110011010"), -- 3.2 + 2.6 = 5.8
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111111010011001100110011001100"), -- 2.6 + -1.8 = 0.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000000011001100110011001101"), -- -0.3 + 2.5 = 2.2
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"00111111010011001100110011001100"), -- 3 + -2.2 = 0.8
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000100000000000000000000000"), -- 0.3 + 3.7 = 4
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000001100110011001100110011"), -- -2.1 + -0.7 = -2.8
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101000110011001100110011"), -- 2.1 + 3 = 5.1
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000001000000000000000000000"), -- -3.5 + 1 = -2.5
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"10111111100011001100110011001110"), -- -3.7 + 2.6 = -1.1
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111110000000000000000000000"), -- 1.5 + -0 = 1.5
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"00111111000000000000000000000000"), -- 1.4 + -0.9 = 0.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111011001100110011001100110"), -- 1.9 + -2.8 = -0.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000000100110011001100110011"), -- 0 + -2.3 = -2.3
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000100010011001100110011010"), -- 1.5 + 2.8 = 4.3
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000101100110011001100110100"), -- 2.2 + 3.4 = 5.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000001100110011001100110011"), -- -0.1 + -2.7 = -2.8
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000000011001100110011001101"), -- -0.6 + -1.6 = -2.2
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000010110011001100110011010"), -- -1.4 + -2 = -3.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111000000000000000000000000"), -- 3 + -2.5 = 0.5
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000100000000000000000000000"), -- -3.8 + -0.2 = -4
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"00111111000110011001100110011000"), -- 2.1 + -1.5 = 0.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000100001100110011001100110"), -- 3.5 + 0.7 = 4.2
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110111001100110011001100"), -- 3.3 + 3.6 = 6.9
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000100000000000000000000000"), -- -3.6 + -0.4 = -4
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000000110011001100110011010"), -- 1.1 + 1.3 = 2.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111101100110011001100110100"), -- 0.3 + 1.1 = 1.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011001100110011001100110"), -- 0.3 + 3.3 = 3.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101110011001100110011010"), -- 3.3 + 2.5 = 5.8
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111111010011001100110011001110"), -- -1.6 + 2.4 = 0.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000000100110011001100110011"), -- 1.4 + 0.9 = 2.3
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"), -- 1.4 + -1.4 = 0
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000011001100110011001100"), -- 0.1 + 2.1 = 2.2
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"10111111110110011001100110011001"), -- -3.1 + 1.4 = -1.7
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111111111001100110011001100110"), -- 2.1 + -0.3 = 1.8
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000100011001100110011001101"), -- 0.8 + 3.6 = 4.4
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000011110011001100110011010"), -- -3.5 + -0.4 = -3.9
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000011001100110011001100110"), -- -2.5 + -1.1 = -3.6
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001110011001100110011001"), -- 3.1 + -0.2 = 2.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"00111111010011001100110011001100"), -- 3 + -2.2 = 0.8
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"10111110100110011001100110100000"), -- 2.1 + -2.4 = -0.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000000010000000000000000000000"), -- -3.6 + 0.6 = -3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000010011001100110011001100"), -- 0.9 + 2.3 = 3.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111110010011001100110011001100"), -- -0.9 + 0.7 = -0.2
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000001100110011001100110011"), -- -1 + -1.8 = -2.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000010000000000000000000000"), -- 0 + 3 = 3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111000000000000000000000000"), -- -0.2 + -0.3 = -0.5
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100100000000000000000000"), -- 1.4 + 3.1 = 4.5
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000110110011001100110011010"), -- -3.4 + -3.4 = -6.8
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000101000110011001100110011"), -- -3.8 + -1.3 = -5.1
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000001110011001100110011010"), -- 0.3 + -3.2 = -2.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000011001100110011001100110"), -- -0.3 + -3.3 = -3.6
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111110010011001100110011001100"), -- -0.6 + 0.8 = 0.2
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000010011001100110011001101"), -- 3.4 + -0.2 = 3.2
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111100000000000000000000001"), -- 2.9 + -1.9 = 1
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"00111111100110011001100110011010"), -- -2.5 + 3.7 = 1.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001000000000000000000000"), -- -0.2 + 2.7 = 2.5
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000101001100110011001100110"), -- 2.4 + 2.8 = 5.2
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000101000000000000000000000"), -- 1.4 + 3.6 = 5
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"10111111011001100110011001101000"), -- 1.3 + -2.2 = -0.9
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111010011001100110011001100"), -- 1.4 + -0.6 = 0.8
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000000010011001100110011001101"), -- -3.3 + 0.1 = -3.2
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000011000000000000000000000"), -- 1.4 + 2.1 = 3.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111111100110011001100110011"), -- 1.9 + -0 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000001100110011001100110"), -- 0 + 2.1 = 2.1
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000110000000000000000000000"), -- -3.3 + -2.7 = -6
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000010110011001100110011010"), -- -0.5 + -2.9 = -3.4
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111000110011001100110011010"), -- 1.2 + -0.6 = 0.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111111010011001100110011001101"), -- 1.5 + -0.7 = 0.8
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000100111001100110011001101"), -- -2.4 + -2.5 = -4.9
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000111011001100110011001101"), -- -3.9 + -3.5 = -7.4
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000100001100110011001100110"), -- -3.6 + -0.6 = -4.2
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000001000000000000000000000"), -- -0.8 + 3.3 = 2.5
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011001100110011001100111"), -- 0.3 + -3.9 = -3.6
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000000110011001100110011010"), -- 2.4 + -0 = 2.4
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000010110011001100110011001"), -- 0.4 + -3.8 = -3.4
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111101111111111111111111111"), -- 1.1 + -2.6 = -1.5
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"10111111110110011001100110011010"), -- -3.8 + 2.1 = -1.7
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000101001100110011001100110"), -- -3.2 + -2 = -5.2
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000001011001100110011001101"), -- 0.3 + 2.4 = 2.7
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000100100110011001100110011"), -- -1.5 + -3.1 = -4.6
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111110010011001100110011001000"), -- -1.9 + 2.1 = 0.2
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000011011001100110011001101"), -- -3.3 + -0.4 = -3.7
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111100011001100110011001100"), -- 1.5 + -2.6 = -1.1
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"00111111111100110011001100110100"), -- -1.5 + 3.4 = 1.9
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000000100110011001100110100"), -- 0.9 + -3.2 = -2.3
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111000000000000000000000010"), -- 2.4 + -1.9 = 0.5
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111110010011001100110011001000"), -- -1.2 + 1.4 = 0.2
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000110100110011001100110011"), -- -3.6 + -3 = -6.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000000100000000000000000000000"), -- 3.5 + 0.5 = 4
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"00111111101100110011001100110100"), -- 2.9 + -1.5 = 1.4
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000000110011001100110011010"), -- 1.8 + 0.6 = 2.4
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101111001100110011001101"), -- 3.7 + 2.2 = 5.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000000000000000000000000"), -- -0.3 + 2.3 = 2
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000101101100110011001100110"), -- 3.6 + 2.1 = 5.7
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111000000000000000000000000"), -- 2.4 + -2.9 = -0.5
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111111001100110011001100111"), -- -1.2 + -0.6 = -1.8
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000010011001100110011001101"), -- 0.8 + 2.4 = 3.2
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111111111100110011001100110100"), -- -0.8 + 2.7 = 1.9
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000010001100110011001100110"), -- -1.7 + -1.4 = -3.1
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"00111111011001100110011001100100"), -- 2.6 + -1.7 = 0.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111110000000000000000000000"), -- -0.9 + -0.6 = -1.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000110110011001100110011010"), -- 3.5 + 3.3 = 6.8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111100110011001100110011000"), -- 3.6 + -2.4 = 1.2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111110100110011001100110011010"), -- 0.2 + -0.5 = -0.3
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101100000000000000000000"), -- -3.9 + -1.6 = -5.5
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000010001100110011001100111"), -- -2.9 + -0.2 = -3.1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001000000000000000000000"), -- 2.5 + -0 = 2.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000000011001100110011001101"), -- 1.9 + 0.3 = 2.2
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000000001100110011001100110"), -- 1.5 + 0.6 = 2.1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000001011001100110011001101"), -- -0.7 + 3.4 = 2.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000000000000000000000000000"), -- 1.1 + 0.9 = 2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111101110011001100110011010000"), -- 2 + -1.9 = 0.1
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111010011001100110011001110"), -- -2.4 + 1.6 = -0.8
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101100110011001100110011"), -- -3 + -2.6 = -5.6
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000101101100110011001100110"), -- -2.3 + -3.4 = -5.7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000110111001100110011001101"), -- 3.7 + 3.2 = 6.9
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111111110110011001100110011010"), -- 1.6 + 0.1 = 1.7
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000001001100110011001100110"), -- -0.8 + -1.8 = -2.6
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000001001100110011001100111"), -- -2.9 + 0.3 = -2.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000001110011001100110011010"), -- 0 + -2.9 = -2.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000100111001100110011001101"), -- -3.5 + -1.4 = -4.9
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000010011001100110011001100"), -- 3.1 + 0.1 = 3.2
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000100011001100110011001101"), -- 3.8 + 0.6 = 4.4
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111110011001100110011001100"), -- 1.7 + -3.3 = -1.6
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000010011001100110011001101"), -- -1.6 + -1.6 = -3.2
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00111111010011001100110011001110"), -- 1.2 + -0.4 = 0.8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000111000000000000000000000"), -- 3.6 + 3.4 = 7
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111100011001100110011001100"), -- 3.6 + -2.5 = 1.1
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000010000000000000000000000"), -- 2 + 1 = 3
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"01000000000110011001100110011010"), -- 3.7 + -1.3 = 2.4
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111110100110011001100110011000"), -- -2.3 + 2.6 = 0.3
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111111001100110011001100111"), -- 1.6 + -3.4 = -1.8
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110101100110011001100110"), -- -3.8 + -2.9 = -6.7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000001011001100110011001101"), -- 3.4 + -0.7 = 2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- 0 + 1.9 = 1.9
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"), -- -2.8 + 2.8 = 0
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"10111111011111111111111111111110"), -- 1.1 + -2.1 = -1
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000101100110011001100110100"), -- -2.7 + -2.9 = -5.6
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000101100000000000000000000"), -- 1.8 + 3.7 = 5.5
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111110110011001100110011001100"), -- 1.5 + -1.1 = 0.4
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111111100011001100110011001101"), -- 0.9 + -2 = -1.1
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000100000110011001100110011"), -- -1.1 + -3 = -4.1
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000100111001100110011001101"), -- -1.7 + -3.2 = -4.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000001000000000000000000000"), -- -3.5 + 1 = -2.5
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000011110011001100110011001"), -- -3.6 + -0.3 = -3.9
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000110100000000000000000000"), -- 3.9 + 2.6 = 6.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111011001100110011001100110"), -- 1.9 + -1 = 0.9
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000101100000000000000000000"), -- -2.1 + -3.4 = -5.5
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000011110011001100110011010"), -- 1.6 + 2.3 = 3.9
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000010110011001100110011010"), -- -1.1 + -2.3 = -3.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000101010011001100110011010"), -- 3 + 2.3 = 5.3
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111111000000000000000000000000"), -- 2.3 + -1.8 = 0.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111101001100110011001100110"), -- 0 + 1.3 = 1.3
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"11000000000001100110011001100110"), -- -3.8 + 1.7 = -2.1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000000110011001100110011010"), -- -0.8 + 3.2 = 2.4
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"10111111100110011001100110011001"), -- -2.6 + 1.4 = -1.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111010011001100110011001101"), -- -0.6 + -0.2 = -0.8
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000110111001100110011001101"), -- 3.4 + 3.5 = 6.9
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000000100110011001100110011"), -- 2.3 + -0 = 2.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111000000000000000000000000"), -- -0.2 + 0.7 = 0.5
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111100110011001100110011001"), -- -3.1 + 1.9 = -1.2
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111001100110011001100110010"), -- -2.3 + 1.6 = -0.7
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000100100000000000000000000"), -- -1.1 + -3.4 = -4.5
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111101001100110011001100111"), -- -2.9 + 1.6 = -1.3
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100101100110011001100110"), -- 1.6 + 3.1 = 4.7
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000011001100110011001100110"), -- -1.8 + -1.8 = -3.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"00111111101001100110011001100111"), -- 2.7 + -1.4 = 1.3
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111110010011001100110011010000"), -- 2.5 + -2.7 = -0.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000100001100110011001100110"), -- 2.8 + 1.4 = 4.2
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000010011001100110011001101"), -- -3.2 + -0 = -3.2
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101000000000000000000000"), -- -3.4 + -1.6 = -5
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000000110011001100110011010"), -- 0.6 + 1.8 = 2.4
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111111110000000000000000000001"), -- -2.4 + 0.9 = -1.5
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111111000000000000000000000000"), -- 1.7 + -1.2 = 0.5
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111110100110011001100110011100"), -- -0.9 + 1.2 = 0.3
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000001000000000000000000000"), -- 0.8 + -3.3 = -2.5
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"00111111000110011001100110011100"), -- 3.7 + -3.1 = 0.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000001001100110011001100111"), -- -1.3 + 3.9 = 2.6
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001011001100110011001101"), -- 2.9 + -0.2 = 2.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000101110011001100110011010"), -- -3.6 + -2.2 = -5.8
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000110101100110011001100110"), -- -2.9 + -3.8 = -6.7
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111011001100110011001100100"), -- -2.1 + 1.2 = -0.9
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000010000000000000000000000"), -- 3.1 + -0.1 = 3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"10111111110000000000000000000000"), -- -2.5 + 1 = -1.5
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001001100110011001100110"), -- 2.6 + -0 = 2.6
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111110010011001100110011001110"), -- 0.4 + -0.6 = -0.2
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111111001100110011001100111"), -- -2.4 + 0.6 = -1.8
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000000100110011001100110011"), -- 0.2 + -2.5 = -2.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000100011001100110011001101"), -- -3.5 + -0.9 = -4.4
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000010100110011001100110100"), -- -0.9 + -2.4 = -3.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111111110110011001100110011010"), -- -3.5 + 1.8 = -1.7
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000011100110011001100110100"), -- -1.6 + -2.2 = -3.8
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000110010011001100110011010"), -- -3.3 + -3 = -6.3
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111000110011001100110011010"), -- 0.3 + 0.3 = 0.6
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000010000000000000000000000"), -- 1.7 + 1.3 = 3
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000001100110011001100110011"), -- -3 + 0.2 = -2.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"00111110100110011001100110100000"), -- 3.9 + -3.6 = 0.3
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"10111111100110011001100110011010"), -- 1 + -2.2 = -1.2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111011001100110011001101000"), -- 2 + -2.9 = -0.9
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000100001100110011001100111"), -- -0.8 + -3.4 = -4.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111010011001100110011001101"), -- -0.7 + -0.1 = -0.8
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111110010011001100110011001000"), -- 1.3 + -1.1 = 0.2
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000101010011001100110011010"), -- -3.5 + -1.8 = -5.3
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111110000000000000000000000"), -- -2.3 + 3.8 = 1.5
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111011001100110011001101000"), -- 3 + -3.9 = -0.9
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"00111110010011001100110011010000"), -- 3.9 + -3.7 = 0.2
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00111111100110011001100110011010"), -- -1.3 + 2.5 = 1.2
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"00111111101100110011001100110100"), -- -2.3 + 3.7 = 1.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000100110011001100110011"), -- 0 + 2.3 = 2.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111110000000000000000000001"), -- 3.4 + -1.9 = 1.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000110000000000000000000000"), -- 3.5 + 2.5 = 6
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000110011001100110011001101"), -- 3.2 + 3.2 = 6.4
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"10111110010011001100110011010000"), -- 2 + -2.2 = -0.2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111101100110011001100110100"), -- -0.3 + -1.1 = -1.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000110111001100110011001101"), -- 3 + 3.9 = 6.9
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010001100110011001100110"), -- -0.2 + 3.3 = 3.1
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000001100110011001100110011"), -- 2 + 0.8 = 2.8
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111101110011001100110011001101"), -- -0.1 + 0.2 = 0.1
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111000110011001100110011000"), -- -2.1 + 1.5 = -0.6
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111111110000000000000000000000"), -- 1.4 + 0.1 = 1.5
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111100110011001100110011010"), -- -0.3 + -0.9 = -1.2
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000101000000000000000000000"), -- -2.6 + -2.4 = -5
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111111001100110011001100110100"), -- -3.5 + 2.8 = -0.7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000101110011001100110011010"), -- -2.8 + -3 = -5.8
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101000110011001100110100"), -- 2.9 + 2.2 = 5.1
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111111001100110011001100110"), -- 0.8 + 1 = 1.8
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000010000000000000000000000"), -- 0.5 + 2.5 = 3
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000001110011001100110011001"), -- 0.8 + 2.1 = 2.9
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111111100000000000000000000000"), -- 1.5 + -0.5 = 1
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000101010011001100110011010"), -- -3.8 + -1.5 = -5.3
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111101111111111111111111111"), -- -3.1 + 1.6 = -1.5
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111110110011001100110011001100"), -- 1.5 + -1.9 = -0.4
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000000000000000000000000000"), -- 1.2 + 0.8 = 2
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000100010011001100110011010"), -- 2.7 + 1.6 = 4.3
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000001000000000000000000000"), -- 1.7 + 0.8 = 2.5
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000011011001100110011001101"), -- 0.2 + -3.9 = -3.7
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111111101001100110011001100110"), -- 1 + -2.3 = -1.3
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000101010011001100110011010"), -- 3.3 + 2 = 5.3
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000011000000000000000000000"), -- -2.7 + -0.8 = -3.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111000110011001100110011000"), -- -3.2 + 3.8 = 0.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- 0 + 3.2 = 3.2
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111100110011001100110011010"), -- -3.2 + 2 = -1.2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111110011001100110011001100"), -- 0.7 + 0.9 = 1.6
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111111101100110011001100110011"), -- 1.9 + -0.5 = 1.4
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111111011111111111111111111111"), -- 1.8 + -0.8 = 1
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000100100000000000000000000"), -- -3.8 + -0.7 = -4.5
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000100100110011001100110011"), -- 1.3 + 3.3 = 4.6
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111111001100110011001100110100"), -- -1.1 + 0.4 = -0.7
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000100010011001100110011010"), -- -0.6 + -3.7 = -4.3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111111010011001100110011001100"), -- -0.5 + 1.3 = 0.8
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111110010011001100110011001000"), -- -1.4 + 1.2 = -0.2
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000110100000000000000000000"), -- -3.1 + -3.4 = -6.5
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111111100000000000000000000000"), -- -2.6 + 3.6 = 1
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000101001100110011001100110"), -- 1.4 + 3.8 = 5.2
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111101001100110011001100110"), -- 1.5 + -2.8 = -1.3
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111100000000000000000000000"), -- 2.3 + -3.3 = -1
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000110000000000000000000000"), -- 3.1 + 2.9 = 6
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000000001100110011001100110"), -- 1.9 + 0.2 = 2.1
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000010011001100110011001101"), -- -3.9 + 0.7 = -3.2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"00111111000000000000000000000000"), -- -2.5 + 3 = 0.5
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111111011001100110011001101000"), -- -2 + 2.9 = 0.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"00111111100110011001100110011001"), -- 2.8 + -1.6 = 1.2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111111100011001100110011001100"), -- 2 + -3.1 = -1.1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000100000000000000000000000"), -- -0.7 + -3.3 = -4
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111100011001100110011001101"), -- 1.1 + -0 = 1.1
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000011000000000000000000000"), -- 3.4 + 0.1 = 3.5
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000010100110011001100110100"), -- -2.2 + -1.1 = -3.3
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"00111111101001100110011001100110"), -- 3 + -1.7 = 1.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000001000000000000000000000"), -- 0.6 + 1.9 = 2.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000001001100110011001100110"), -- 0 + 2.6 = 2.6
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111101110011001100110011000000"), -- 2.1 + -2 = 0.0999999
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000101111001100110011001101"), -- -3.7 + -2.2 = -5.9
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000001011001100110011001101"), -- 1.2 + 1.5 = 2.7
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000000000000000000000000000"), -- -1.3 + 3.3 = 2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000101000110011001100110100"), -- 2.4 + 2.7 = 5.1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000100100110011001100110011"), -- -0.8 + -3.8 = -4.6
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000010011001100110011001100"), -- -0.6 + -2.6 = -3.2
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000111010011001100110011010"), -- -3.5 + -3.8 = -7.3
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000010000000000000000000000"), -- 0.4 + 2.6 = 3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111100110011001100110011010"), -- 2.6 + -3.8 = -1.2
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000100010011001100110011010"), -- 0.9 + 3.4 = 4.3
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"00111111001100110011001100110100"), -- -2.7 + 3.4 = 0.7
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"10111111101100110011001100110100"), -- -3.5 + 2.1 = -1.4
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111110010011001100110011000000"), -- 2.6 + -2.4 = 0.2
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"10111111100000000000000000000000"), -- 2.5 + -3.5 = -1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000000011001100110011001100"), -- 0.6 + -2.8 = -2.2
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000010001100110011001100110"), -- -1.9 + -1.2 = -3.1
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000000100110011001100110011"), -- -2.7 + 0.4 = -2.3
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000100000110011001100110100"), -- -2.9 + -1.2 = -4.1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"), -- 2.5 + -2.5 = 0
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111111001100110011001100110"), -- 1.8 + -0 = 1.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111001100110011001100110100"), -- -0.3 + -0.4 = -0.7
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000001000000000000000000000"), -- 2.3 + 0.2 = 2.5
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000101111001100110011001100"), -- -2.8 + -3.1 = -5.9
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111101110011001100110011000000"), -- 2.6 + -2.5 = 0.0999999
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000100101100110011001100110"), -- -2.7 + -2 = -4.7
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110000000000000000000000"), -- 2.4 + 3.6 = 6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111111100000000000000000000000"), -- 1.5 + -0.5 = 1
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000000001100110011001100110"), -- 0.7 + 1.4 = 2.1
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000001100110011001100110011"), -- 2 + 0.8 = 2.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000110100000000000000000000"), -- 3.8 + 2.7 = 6.5
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000001011001100110011001100"), -- 2.6 + 0.1 = 2.7
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100000000000000000000000"), -- 0.9 + 3.1 = 4
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010100110011001100110011"), -- -0.2 + -3.1 = -3.3
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111100000000000000000000000"), -- -0.7 + 1.7 = 1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111111001100110011001100110"), -- -0.8 + 2.6 = 1.8
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111100110011001100110011010"), -- -0.7 + 1.9 = 1.2
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000010100110011001100110011"), -- -2 + -1.3 = -3.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000101100110011001100110011"), -- -3.6 + -2 = -5.6
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000100110011001100110011010"), -- 2.9 + 1.9 = 4.8
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"10111101110011001100110011000000"), -- -3.3 + 3.2 = -0.0999999
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"00111110100110011001100110011000"), -- -3.4 + 3.7 = 0.3
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000100000110011001100110011"), -- -1.5 + -2.6 = -4.1
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"), -- 1.1 + -1.1 = 0
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111100000000000000000000000"), -- -3 + 2 = -1
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000110100000000000000000000"), -- 3.7 + 2.8 = 6.5
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"00111111101100110011001100110100"), -- -2 + 3.4 = 1.4
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000100000000000000000000000"), -- 1.9 + 2.1 = 4
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111000000000000000000000000"), -- 0.1 + 0.4 = 0.5
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000001110011001100110011010"), -- 0.5 + -3.4 = -2.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000000011001100110011001101"), -- -0.3 + -1.9 = -2.2
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111111001100110011001100110"), -- 0.9 + 0.9 = 1.8
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"00111111000000000000000000000000"), -- 3.3 + -2.8 = 0.5
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000011000000000000000000000"), -- 2.7 + 0.8 = 3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- 0 + 3.2 = 3.2
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110000000000000000000000"), -- -3.1 + -2.9 = -6
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111100110011001100110011010"), -- -0.7 + 1.9 = 1.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111000000000000000000000001"), -- -0.7 + 1.2 = 0.5
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000101000110011001100110011"), -- 3.7 + 1.4 = 5.1
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000110000000000000000000000"), -- 3.1 + 2.9 = 6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000001011001100110011001101"), -- 1.5 + 1.2 = 2.7
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111010011001100110011001100"), -- -2 + 2.8 = 0.8
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000010100110011001100110011"), -- 3.3 + -0 = 3.3
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000100110011001100110011010"), -- -1.5 + -3.3 = -4.8
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111110110011001100110011010000"), -- -2.3 + 2.7 = 0.4
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111000110011001100110011000"), -- 3.1 + -2.5 = 0.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111100000000000000000000000"), -- -1.3 + 2.3 = 1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000000001100110011001100110"), -- 2.5 + -0.4 = 2.1
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000011100110011001100110100"), -- 1.1 + 2.7 = 3.8
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000010110011001100110011010"), -- 1.8 + 1.6 = 3.4
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000011100110011001100110011"), -- -2.5 + -1.3 = -3.8
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000011100110011001100110011"), -- -3.8 + -0 = -3.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000000000000000000000000000"), -- -0.3 + -1.7 = -2
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000011110011001100110011001"), -- 2.1 + 1.8 = 3.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000111000000000000000000000"), -- -3.5 + -3.5 = -7
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111110110011001100110011010000"), -- -2.5 + 2.9 = 0.4
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111111001100110011001100111"), -- 1.1 + -2.9 = -1.8
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111111000110011001100110011010"), -- -0.8 + 0.2 = -0.6
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000001001100110011001100111"), -- 0.4 + 2.2 = 2.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000000000000000000000000000000"), -- 1.5 + 0.5 = 2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000000001100110011001100110"), -- 2.8 + -0.7 = 2.1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"00111111100110011001100110011001"), -- 2.1 + -0.9 = 1.2
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000110000000000000000000000"), -- 2.7 + 3.3 = 6
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000100000110011001100110011"), -- -0.3 + -3.8 = -4.1
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000100000000000000000000000"), -- -3.7 + -0.3 = -4
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"10111111100000000000000000000001"), -- 1.4 + -2.4 = -1
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000101100110011001100110100"), -- 1.7 + 3.9 = 5.6
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000010110011001100110011010"), -- 2.2 + 1.2 = 3.4
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111111001100110011001100110"), -- -3 + 1.2 = -1.8
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000001011001100110011001101"), -- 0.5 + 2.2 = 2.7
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"00111111001100110011001100110100"), -- -2.3 + 3 = 0.7
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000100000000000000000000000"), -- 0.3 + 3.7 = 4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111111111100110011001100110100"), -- 2.7 + -0.8 = 1.9
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000000110011001100110011001"), -- -1.2 + 3.6 = 2.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"10111111000000000000000000000000"), -- 3 + -3.5 = -0.5
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111101111111111111111111111"), -- -3.1 + 1.6 = -1.5
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000101101100110011001100110"), -- -3.8 + -1.9 = -5.7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000000000000000000000000000"), -- 3.7 + -1.7 = 2
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000100110011001100110011010"), -- -2.1 + -2.7 = -4.8
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000110101100110011001100110"), -- 2.8 + 3.9 = 6.7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111100011001100110011001110"), -- -2.8 + 3.9 = 1.1
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000001100110011001100110100"), -- -2.4 + -0.4 = -2.8
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000010110011001100110011010"), -- 2.4 + 1 = 3.4
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00111111111001100110011001100111"), -- 2.2 + -0.4 = 1.8
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111110010011001100110011001100"), -- 0.5 + -0.3 = 0.2
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111010011001100110011001100"), -- -2 + 2.8 = 0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011011001100110011001101"), -- 0 + 3.7 = 3.7
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"00111111100110011001100110011010"), -- -2 + 3.2 = 1.2
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"10111111110000000000000000000000"), -- -3.8 + 2.3 = -1.5
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000101000110011001100110100"), -- -1.7 + -3.4 = -5.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"00111101110011001100110011000000"), -- -1.2 + 1.3 = 0.0999999
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111111100110011001100110010"), -- 0.7 + -2.6 = -1.9
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000110101100110011001100110"), -- -3 + -3.7 = -6.7
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00111111110011001100110011001101"), -- 2 + -0.4 = 1.6
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111110110011001100110011010000"), -- 1.3 + -1.7 = -0.4
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000000000000000000000000000"), -- -2.7 + 0.7 = -2
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111110011001100110011001100"), -- 1 + -2.6 = -1.6
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000011011001100110011001101"), -- -3.9 + 0.2 = -3.7
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111110000000000000000000000"), -- 1.6 + -0.1 = 1.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- 0 + 3.2 = 3.2
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"10111111000110011001100110011000"), -- -2.3 + 1.7 = -0.6
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000010110011001100110011001"), -- -3.6 + 0.2 = -3.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111110010011001100110011010000"), -- -1.1 + 0.9 = -0.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111101001100110011001100111"), -- 3.2 + -1.9 = 1.3
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000110100000000000000000000"), -- -3 + -3.5 = -6.5
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000100100110011001100110100"), -- 2.9 + 1.7 = 4.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000100110011001100110100"), -- -0.1 + 2.4 = 2.3
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111100011001100110011001100"), -- -2.2 + 3.3 = 1.1
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111011001100110011001101000"), -- -3 + 3.9 = 0.9
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000100011001100110011001101"), -- -2.8 + -1.6 = -4.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000100100110011001100110011"), -- -1.1 + -3.5 = -4.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111110110011001100110011001100"), -- -1.3 + 0.9 = -0.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000001110011001100110011001"), -- -3.3 + 0.4 = -2.9
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000100011001100110011001101"), -- 3.2 + 1.2 = 4.4
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111101100110011001100110011"), -- 3.3 + -1.9 = 1.4
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000001110011001100110011010"), -- -2.4 + -0.5 = -2.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000001001100110011001100110"), -- -0.9 + -1.7 = -2.6
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000001100110011001100110011"), -- 3.1 + -0.3 = 2.8
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111101001100110011001100111"), -- -0.9 + 2.2 = 1.3
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"10111111010011001100110011001101"), -- -0.1 + -0.7 = -0.8
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000011011001100110011001100"), -- 2.8 + 0.9 = 3.7
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000101100110011001100110100"), -- -3.4 + -2.2 = -5.6
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111110110011001100110011001110"), -- -0.8 + 1.2 = 0.4
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000100000000000000000000000"), -- 2.9 + 1.1 = 4
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000101001100110011001100110"), -- 2.8 + 2.4 = 5.2
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000010011001100110011001101"), -- -3.2 + -0 = -3.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111111001100110011001100110"), -- -0.5 + 2.3 = 1.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000101110011001100110011010"), -- 3.8 + 2 = 5.8
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111111010011001100110011001101"), -- -1.5 + 0.7 = -0.8
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000000000000000000000000000"), -- -1.2 + 3.2 = 2
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000100010011001100110011010"), -- -0.8 + -3.5 = -4.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"10111111101100110011001100110010"), -- -3.6 + 2.2 = -1.4
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000000001100110011001100110"), -- 1.4 + -3.5 = -2.1
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000001100110011001100110011"), -- -1.3 + -1.5 = -2.8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000000100000110011001100110011"), -- 3.6 + 0.5 = 4.1
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000100001100110011001100110"), -- 3.8 + 0.4 = 4.2
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"10111111101100110011001100110100"), -- 1.8 + -3.2 = -1.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000100001100110011001100110"), -- -3.3 + -0.9 = -4.2
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000000011001100110011001101"), -- 1 + 1.2 = 2.2
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000000110011001100110011001"), -- -2.8 + 0.4 = -2.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111110110011001100110011001101"), -- 0 + -0.4 = -0.4
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000100011001100110011001101"), -- 2.9 + 1.5 = 4.4
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000000110011001100110011010"), -- 2.5 + -0.1 = 2.4
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"10111111111001100110011001100110"), -- -3.5 + 1.7 = -1.8
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111111100000000000000000000000"), -- -3.5 + 2.5 = -1
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000001110011001100110011010"), -- 0.1 + -3 = -2.9
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000101000000000000000000000"), -- 3.3 + 1.7 = 5
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000100101100110011001100110"), -- 2.1 + 2.6 = 4.7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111001100110011001100110100"), -- -2.8 + 3.5 = 0.7
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000001100110011001100111"), -- 0.3 + -2.4 = -2.1
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101110011001100110011010"), -- -3.2 + -2.6 = -5.8
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111101110011001100110011100000"), -- -2.3 + 2.4 = 0.1
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"11000000000100110011001100110100"), -- -3.4 + 1.1 = -2.3
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"01000000000011001100110011001101"), -- 3.5 + -1.3 = 2.2
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000100001100110011001100110"), -- 2.1 + 2.1 = 4.2
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000010001100110011001100110"), -- 0.6 + -3.7 = -3.1
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111100110011001100110011"), -- 0.1 + 1.8 = 1.9
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000010110011001100110011010"), -- 0.5 + 2.9 = 3.4
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111101001100110011001101000"), -- 3.4 + -2.1 = 1.3
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000100000110011001100110011"), -- -0.7 + -3.4 = -4.1
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000000000000000000000000"), -- -0.3 + 2.3 = 2
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111100110011001100110011010"), -- -2.6 + 3.8 = 1.2
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000101000110011001100110011"), -- -3.7 + -1.4 = -5.1
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"10111111111100110011001100110011"), -- -0.4 + -1.5 = -1.9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111111110110011001100110011010"), -- 2.9 + -1.2 = 1.7
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000001000000000000000000000"), -- 1.5 + 1 = 2.5
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000000001011001100110011001101"), -- 2.2 + 0.5 = 2.7
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"00111111001100110011001100110100"), -- 2 + -1.3 = 0.7
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111110010011001100110011010000"), -- 1.4 + -1.6 = -0.2
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000101011001100110011001100"), -- -2.6 + -2.8 = -5.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"10111101110011001100110011000000"), -- -1.8 + 1.7 = -0.0999999
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111010011001100110011001101"), -- 0 + 0.8 = 0.8
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000100110011001100110011010"), -- 2.6 + 2.2 = 4.8
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000000011001100110011001100"), -- -1.6 + 3.8 = 2.2
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111111000110011001100110011100"), -- 2.1 + -2.7 = -0.6
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111110110011001100110011001100"), -- -1.9 + 2.3 = 0.4
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000011100110011001100110011"), -- 1.2 + 2.6 = 3.8
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111010011001100110011001110"), -- 2.7 + -1.9 = 0.8
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111100000000000000000000000"), -- -0.2 + 1.2 = 1
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000101100000000000000000000"), -- -2.2 + -3.3 = -5.5
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000000110011001100110011010"), -- 1.1 + -3.5 = -2.4
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"10111111001100110011001100110100"), -- 1.7 + -2.4 = -0.7
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000100011001100110011001101"), -- -0.5 + -3.9 = -4.4
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"00111110100110011001100110011000"), -- 2.6 + -2.3 = 0.3
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111100110011001100110011001"), -- 1.8 + -0.6 = 1.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000101010011001100110011010"), -- 2.8 + 2.5 = 5.3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000011000000000000000000000"), -- 2.6 + 0.9 = 3.5
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000100110011001100110011010"), -- 1.1 + 3.7 = 4.8
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"10111111111100110011001100110010"), -- -3.6 + 1.7 = -1.9
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000000100110011001100110011"), -- -1 + 3.3 = 2.3
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000100101100110011001100110"), -- -2 + -2.7 = -4.7
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"00111110110011001100110011010000"), -- 1.7 + -1.3 = 0.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000100001100110011001100111"), -- 0.3 + 3.9 = 4.2
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000010011001100110011001101"), -- -2.4 + -0.8 = -3.2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000100101100110011001100110"), -- 2 + 2.7 = 4.7
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000010001100110011001100111"), -- 0.1 + -3.2 = -3.1
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000010000000000000000000000"), -- -2.8 + -0.2 = -3
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000101111001100110011001101"), -- -3 + -2.9 = -5.9
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"00111111001100110011001100110100"), -- 3.7 + -3 = 0.7
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000000110011001100110011010"), -- 1.5 + -3.9 = -2.4
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111001100110011001100110011"), -- 0.8 + -0.1 = 0.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000010001100110011001100110"), -- -3.6 + 0.5 = -3.1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000010001100110011001100110"), -- -0.8 + -2.3 = -3.1
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111000000000000000000000000"), -- -1.1 + 1.6 = 0.5
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000001011001100110011001101"), -- -1.2 + 3.9 = 2.7
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111111100110011001100110100"), -- -3.4 + 1.5 = -1.9
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00111111111100110011001100110010"), -- -1.2 + 3.1 = 1.9
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110000000000000000000000"), -- -3.1 + -2.9 = -6
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000100001100110011001100110"), -- -0.9 + -3.3 = -4.2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101011001100110011001101"), -- 2.4 + 3 = 5.4
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000101101100110011001100110"), -- 2 + 3.7 = 5.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000101100000000000000000000"), -- 2.2 + 3.3 = 5.5
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111101001100110011001100110"), -- 0.6 + 0.7 = 1.3
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111000000000000000000000000"), -- 1.5 + -1 = 0.5
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"00111111011001100110011001100100"), -- 2.6 + -1.7 = 0.9
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000000001100110011001100110"), -- 0.6 + 1.5 = 2.1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000010011001100110011001101"), -- -0.7 + 3.9 = 3.2
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000100000110011001100110011"), -- 3.9 + 0.2 = 4.1
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000100001100110011001100110"), -- -1.9 + -2.3 = -4.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000100111001100110011001101"), -- 3.2 + 1.7 = 4.9
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000100011001100110011001101"), -- -1.2 + -3.2 = -4.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000010110011001100110011010"), -- -1.8 + -1.6 = -3.4
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000011011001100110011001100"), -- 2.6 + 1.1 = 3.7
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000011011001100110011001101"), -- 3.5 + 0.2 = 3.7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000100010011001100110011010"), -- 3.4 + 0.9 = 4.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111000000000000000000000000"), -- -0.2 + 0.7 = 0.5
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010110011001100110011010"), -- 0.2 + 3.2 = 3.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111111100110011001100110100"), -- 0.3 + 1.6 = 1.9
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"10111111000110011001100110011100"), -- -3.9 + 3.3 = -0.6
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000011011001100110011001100"), -- 2.3 + 1.4 = 3.7
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000001110011001100110011010"), -- 0.6 + -3.5 = -2.9
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111111101100110011001100110100"), -- -2.2 + 0.8 = -1.4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000100110011001100110011010"), -- 2.7 + 2.1 = 4.8
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000011011001100110011001101"), -- -3.7 + -0 = -3.7
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000011100110011001100110011"), -- -3.3 + -0.5 = -3.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111110110011001100110011001100"), -- 1.4 + -1.8 = -0.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000111000110011001100110100"), -- -3.7 + -3.4 = -7.1
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000000001100110011001100110"), -- 0.9 + -3 = -2.1
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111111110110011001100110011010"), -- -2.4 + 0.7 = -1.7
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111100011001100110011001101"), -- 0.5 + -1.6 = -1.1
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000010100110011001100110011"), -- 3.5 + -0.2 = 3.3
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000110001100110011001100110"), -- 3.9 + 2.3 = 6.2
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000000011001100110011001101"), -- -3.4 + 1.2 = -2.2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000101100110011001100110011"), -- -2.5 + -3.1 = -5.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000100010011001100110011010"), -- 2 + 2.3 = 4.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111111110110011001100110011010"), -- -1.2 + 2.9 = 1.7
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000011011001100110011001101"), -- 2.7 + 1 = 3.7
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"10111101110011001100110011000000"), -- -3.1 + 3 = -0.0999999
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"00111111001100110011001100110011"), -- -0.7 + 1.4 = 0.7
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111000000000000000000000000"), -- 3.3 + -3.8 = -0.5
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"00111111011001100110011001100110"), -- 1.8 + -0.9 = 0.9
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000100001100110011001100110"), -- -1.9 + -2.3 = -4.2
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000100100000000000000000000"), -- 3.3 + 1.2 = 4.5
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000011110011001100110011010"), -- 2.2 + 1.7 = 3.9
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000100001100110011001100110"), -- 1.6 + 2.6 = 4.2
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111110010011001100110011001110"), -- -0.1 + 0.3 = 0.2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111110100110011001100110011010"), -- -0.3 + 0.6 = 0.3
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000101011001100110011001100"), -- -3.3 + -2.1 = -5.4
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000000000000000000000000000"), -- 0.1 + 1.9 = 2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000001110011001100110011010"), -- -0.9 + 3.8 = 2.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111111100110011001100110011"), -- -0.9 + 2.8 = 1.9
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000101000000000000000000000"), -- -2 + -3 = -5
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111111000110011001100110011010"), -- -1.5 + 0.9 = -0.6
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"00111111110110011001100110011010"), -- 1 + 0.7 = 1.7
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000011011001100110011001101"), -- -0.2 + -3.5 = -3.7
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00111111110000000000000000000000"), -- 1.9 + -0.4 = 1.5
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111001100110011001100110100"), -- -2.7 + 2 = -0.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000101100000000000000000000"), -- 2.2 + 3.3 = 5.5
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000100010011001100110011010"), -- -3.3 + -1 = -4.3
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000010100110011001100110011"), -- -0.3 + 3.6 = 3.3
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"11000000010000000000000000000000"), -- -2.9 + -0.1 = -3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111110110011001100110011010"), -- -0.5 + -1.2 = -1.7
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000000100110011001100110011"), -- 1.3 + -3.6 = -2.3
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000111000000000000000000000"), -- 3.2 + 3.8 = 7
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111110100110011001100110011000"), -- 2.3 + -2 = 0.3
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111110111111111111111111111111"), -- -0.9 + 0.4 = -0.5
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000010110011001100110011010"), -- 0.7 + 2.7 = 3.4
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000110100000000000000000000"), -- 2.6 + 3.9 = 6.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"10111111000000000000000000000000"), -- 2.5 + -3 = -0.5
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111000000000000000000000000"), -- -1.3 + 1.8 = 0.5
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111001100110011001100110100"), -- 2.6 + -3.3 = -0.7
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111101111111111111111111111"), -- 2.1 + -0.6 = 1.5
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000001000000000000000000000"), -- 1.6 + 0.9 = 2.5
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000100100000000000000000000"), -- -3.8 + -0.7 = -4.5
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111111011111111111111111111111"), -- -1.3 + 0.3 = -1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000101010011001100110011010"), -- 2.1 + 3.2 = 5.3
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111101100110011001100110010"), -- 2.2 + -3.6 = -1.4
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00111111110011001100110011001101"), -- -0.9 + 2.5 = 1.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"10111111101100110011001100110011"), -- -0.1 + -1.3 = -1.4
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000100000000000000000000000"), -- -3.2 + -0.8 = -4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"10111110110011001100110011001000"), -- -3.8 + 3.4 = -0.4
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111101001100110011001100110"), -- -0.7 + -0.6 = -1.3
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000011001100110011001100110"), -- -1.9 + -1.7 = -3.6
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000000100110011001100110100"), -- 0.6 + 1.7 = 2.3
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000100000000000000000000000"), -- -3.8 + -0.2 = -4
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000001100110011001100110011"), -- -0.4 + 3.2 = 2.8
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000001000000000000000000000"), -- 3 + -0.5 = 2.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111111100110011001100110011"), -- 0.4 + 1.5 = 1.9
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000001100110011001100110011"), -- 1 + 1.8 = 2.8
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111101001100110011001100110"), -- 0.6 + -1.9 = -1.3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000000100110011001100110011"), -- 0.9 + 1.4 = 2.3
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000000001100110011001100110"), -- 0.4 + -2.5 = -2.1
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"10111111110011001100110011001100"), -- -2.1 + 0.5 = -1.6
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000100111001100110011001101"), -- 2.4 + 2.5 = 4.9
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111110100110011001100110011010"), -- 0.6 + -0.3 = 0.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000100101100110011001100110"), -- -3.5 + -1.2 = -4.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111001100110011001100110100"), -- 2.6 + -3.3 = -0.7
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111100011001100110011001101"), -- -0.5 + -0.6 = -1.1
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000010001100110011001100110"), -- 1.2 + 1.9 = 3.1
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"00111110010011001100110011010000"), -- 3 + -2.8 = 0.2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"10111101110011001100110011010000"), -- -1.1 + 1 = -0.1
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000110001100110011001100110"), -- -3.5 + -2.7 = -6.2
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000000011001100110011001101"), -- 2.3 + -0.1 = 2.2
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000100010011001100110011010"), -- 1.5 + 2.8 = 4.3
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000100100110011001100110100"), -- 1.2 + 3.4 = 4.6
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"10111111111001100110011001101000"), -- -3.9 + 2.1 = -1.8
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111110110011001100110011001100"), -- 1.2 + -1.6 = -0.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"10111111000110011001100110011000"), -- -3.3 + 2.7 = -0.6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00111111100011001100110011001101"), -- -1.4 + 2.5 = 1.1
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"10111111000000000000000000000010"), -- 1.9 + -2.4 = -0.5
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000010001100110011001100110"), -- 0.8 + 2.3 = 3.1
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000001001100110011001100110"), -- -1.8 + -0.8 = -2.6
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000001100110011001100110011"), -- -1.9 + -0.9 = -2.8
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"10111111100110011001100110011010"), -- -1.5 + 0.3 = -1.2
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111000110011001100110011100"), -- 2.3 + -2.9 = -0.6
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000001000000000000000000000"), -- 3 + -0.5 = 2.5
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000010001100110011001100111"), -- -0.3 + 3.4 = 3.1
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000100011001100110011001101"), -- 3.6 + 0.8 = 4.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000001011001100110011001101"), -- -3.7 + 1 = -2.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111101110011001100110011001101"), -- 0 + -0.1 = -0.1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111010011001100110011001101"), -- -0.8 + -0 = -0.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000000001000000000000000000000"), -- -2.6 + 0.1 = -2.5
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111101110011001100110011000000"), -- -2.7 + 2.8 = 0.0999999
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000010110011001100110011010"), -- 1.2 + 2.2 = 3.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"11000000010110011001100110011001"), -- -3.3 + -0.1 = -3.4
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"00111111110110011001100110011010"), -- -2 + 3.7 = 1.7
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111111100110011001100110100"), -- -0.2 + -1.7 = -1.9
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111111001100110011001100110"), -- 1.5 + 0.3 = 1.8
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000110110011001100110011010"), -- 3.2 + 3.6 = 6.8
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111101100110011001100110100"), -- -2.5 + 3.9 = 1.4
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000110010011001100110011010"), -- -2.5 + -3.8 = -6.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111111111100110011001100110100"), -- -1 + 2.9 = 1.9
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000100101100110011001100111"), -- 3.9 + 0.8 = 4.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111110100110011001100110011100"), -- 2.2 + -1.9 = 0.3
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000100111001100110011001101"), -- -2 + -2.9 = -4.9
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111101110011001100110011010000"), -- -1.8 + 1.9 = 0.1
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000001001100110011001100110"), -- -3.1 + 0.5 = -2.6
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000001100110011001100110011"), -- 0.3 + -3.1 = -2.8
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000101010011001100110011010"), -- 1.8 + 3.5 = 5.3
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111111001100110011001100110"), -- -1.8 + -0 = -1.8
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000110000110011001100110011"), -- 2.3 + 3.8 = 6.1
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000011001100110011001100111"), -- -2.9 + -0.7 = -3.6
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000011001100110011001100110"), -- -2.6 + -1 = -3.6
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111100110011001100110011010"), -- 0 + -1.2 = -1.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000001011001100110011001101"), -- -0.5 + 3.2 = 2.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111000000000000000000000000"), -- 1.1 + -0.6 = 0.5
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000100000110011001100110011"), -- -3.7 + -0.4 = -4.1
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111110110011001100110011001000"), -- 3.2 + -3.6 = -0.4
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000010000000000000000000000"), -- -2.3 + -0.7 = -3
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000001001100110011001100111"), -- -1.3 + 3.9 = 2.6
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"00111111110011001100110011001100"), -- 1.8 + -0.2 = 1.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111111101001100110011001100110"), -- 2 + -0.7 = 1.3
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000101010011001100110011010"), -- -3.1 + -2.2 = -5.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111111111111111111111111111"), -- -3.6 + 1.6 = -2
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111110110011001100110011010"), -- -1.6 + -0.1 = -1.7
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000001110011001100110011010"), -- 2.9 + -0 = 2.9
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111100000000000000000000000"), -- -0.2 + -0.8 = -1
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111110110011001100110011001"), -- 2.3 + -0.6 = 1.7
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000010100110011001100110100"), -- -2.2 + -1.1 = -3.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111001100110011001100110100"), -- 3.4 + -2.7 = 0.7
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"10111111110110011001100110011010"), -- 1.8 + -3.5 = -1.7
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111001100110011001100110"), -- -0.1 + 1.9 = 1.8
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000100100110011001100110011"), -- -2.7 + -1.9 = -4.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111111110000000000000000000000"), -- 2.7 + -1.2 = 1.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111011001100110011001101000"), -- 2.5 + -3.4 = -0.9
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000100000000000000000000000"), -- -0.1 + -3.9 = -4
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000011000000000000000000000"), -- 0.6 + 2.9 = 3.5
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000100000110011001100110011"), -- 3.8 + 0.3 = 4.1
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000001001100110011001100110"), -- -2.8 + 0.2 = -2.6
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111011001100110011001100110"), -- -1.9 + 2.8 = 0.9
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111110110011001100110011010"), -- 1.2 + -2.9 = -1.7
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111110110011001100110011010"), -- 3.8 + -2.1 = 1.7
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000100011001100110011001101"), -- -1.6 + -2.8 = -4.4
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"10111111000000000000000000000000"), -- -1.5 + 1 = -0.5
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101110011001100110011010"), -- 2.8 + 3 = 5.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000011001100110011001100110"), -- -0.3 + -3.3 = -3.6
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000010110011001100110011010"), -- -1 + -2.4 = -3.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000100110011001100110100"), -- -3.7 + 1.4 = -2.3
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111100011001100110011001101"), -- -0.1 + -1 = -1.1
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000001110011001100110011010"), -- -1.5 + -1.4 = -2.9
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111111100110011001100110011010"), -- -3 + 1.8 = -1.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000000001100110011001100110"), -- 3.2 + -1.1 = 2.1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000001110011001100110011010"), -- 0.6 + -3.5 = -2.9
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111101110011001100110011010000"), -- -1.5 + 1.6 = 0.1
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000110010011001100110011010"), -- -3.3 + -3 = -6.3
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000010110011001100110011010"), -- 1.5 + 1.9 = 3.4
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111010011001100110011001100"), -- -1.8 + 2.6 = 0.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"10111111110000000000000000000000"), -- -2.8 + 1.3 = -1.5
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000011100110011001100110100"), -- -0.6 + -3.2 = -3.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"00111110110011001100110011001000"), -- 3.8 + -3.4 = 0.4
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111010011001100110011001100"), -- 3.5 + -2.7 = 0.8
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000101000000000000000000000"), -- -2.6 + -2.4 = -5
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"10111111000000000000000000000000"), -- -1 + 0.5 = -0.5
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000001100110011001100111"), -- -0.1 + 2.2 = 2.1
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000101010011001100110011010"), -- 3 + 2.3 = 5.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000101100000000000000000000"), -- -3.6 + -1.9 = -5.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"10111111101100110011001100110100"), -- -3.2 + 1.8 = -1.4
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000001110011001100110011010"), -- -1.2 + -1.7 = -2.9
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000101100110011001100110011"), -- 3.5 + 2.1 = 5.6
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001110011001100110011010"), -- -0.4 + -2.5 = -2.9
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000011000000000000000000000"), -- 3.5 + -0 = 3.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000011110011001100110011010"), -- 1.9 + 2 = 3.9
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000101111001100110011001100"), -- -2.1 + -3.8 = -5.9
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000111011001100110011001100"), -- -3.8 + -3.6 = -7.4
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000011110011001100110011010"), -- 3.2 + 0.7 = 3.9
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111101110011001100110011100000"), -- 3.6 + -3.7 = -0.1
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000000011001100110011001101"), -- 1.9 + 0.3 = 2.2
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"10111111100110011001100110011001"), -- -2.6 + 1.4 = -1.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000010011001100110011001101"), -- -0.7 + 3.9 = 3.2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000000110011001100110011010"), -- -1.2 + -1.2 = -2.4
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000011110011001100110011010"), -- 3.7 + 0.2 = 3.9
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000110011001100110011001101"), -- 2.7 + 3.7 = 6.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111111001100110011001100110"), -- -3.3 + 1.5 = -1.8
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111111011001100110011001100111"), -- -1.1 + 0.2 = -0.9
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000101101100110011001100110"), -- -3.9 + -1.8 = -5.7
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000100000110011001100110011"), -- 0.4 + 3.7 = 4.1
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"00111110110011001100110011001101"), -- 0.3 + 0.1 = 0.4
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"00111111000110011001100110011100"), -- -2.3 + 2.9 = 0.6
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000010100110011001100110011"), -- -3.8 + 0.5 = -3.3
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100110011001100110011010"), -- 1.3 + 3.5 = 4.8
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"00111111000110011001100110011010"), -- 1.5 + -0.9 = 0.6
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00111111101001100110011001100110"), -- -1.8 + 3.1 = 1.3
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000001100110011001100110011"), -- -0.8 + 3.6 = 2.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111100110011001100110011010"), -- 3.9 + -2.7 = 1.2
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000100101100110011001100111"), -- -3.9 + -0.8 = -4.7
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"00111111100000000000000000000000"), -- 3.6 + -2.6 = 1
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111111101001100110011001100110"), -- 2.4 + -3.7 = -1.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000001011001100110011001100"), -- -0.6 + 3.3 = 2.7
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000001001100110011001100110"), -- -3.3 + 0.7 = -2.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000011110011001100110011010"), -- -2 + -1.9 = -3.9
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000010001100110011001100110"), -- 1.9 + 1.2 = 3.1
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000001110011001100110011010"), -- -1.1 + -1.8 = -2.9
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111010011001100110011001100"), -- -2.5 + 3.3 = 0.8
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111100000000000000000000000"), -- -2.5 + 3.5 = 1
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000000000100110011001100110011"), -- -3.6 + 1.3 = -2.3
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000000001100110011001100110"), -- 1.9 + 0.2 = 2.1
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000001110011001100110011010"), -- 0.5 + -3.4 = -2.9
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000100100000000000000000000"), -- 0.7 + 3.8 = 4.5
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111000000000000000000000000"), -- 0.6 + -1.1 = -0.5
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000001100110011001100110011"), -- 2.7 + 0.1 = 2.8
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100000000000000000000000"), -- 0.1 + -1.1 = -1
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111111111111111111111111111"), -- -3.1 + 1.1 = -2
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000100110011001100110011010"), -- 1.1 + 3.7 = 4.8
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111110011001100110011001101"), -- 1.7 + -0.1 = 1.6
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000001100110011001100110"), -- -3.5 + 1.4 = -2.1
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111111001100110011001100110"), -- 0.8 + -2.6 = -1.8
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000000001100110011001100110"), -- 1.7 + -3.8 = -2.1
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000001000000000000000000000"), -- -2.2 + -0.3 = -2.5
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000110100110011001100110011"), -- 3.1 + 3.5 = 6.6
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"10111111100110011001100110011010"), -- -0.9 + -0.3 = -1.2
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000011001100110011001100110"), -- 0.5 + 3.1 = 3.6
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111110110011001100110011001"), -- -2.8 + 1.1 = -1.7
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111100000000000000000000000"), -- 2.9 + -3.9 = -1
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111100110011001100110011010"), -- 0.4 + 0.8 = 1.2
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"00111110110011001100110011001110"), -- 0.6 + -0.2 = 0.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000110000110011001100110100"), -- -3.7 + -2.4 = -6.1
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"), -- 3 + -3 = 0
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000011001100110011001100110"), -- -2.1 + -1.5 = -3.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000000100110011001100110011"), -- 2 + 0.3 = 2.3
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000000000000000000000000000"), -- -0.4 + 2.4 = 2
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111111001100110011001100111"), -- 0.6 + 1.2 = 1.8
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"10111111100000000000000000000000"), -- -1.4 + 0.4 = -1
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101100000000000000000000"), -- -3.9 + -1.6 = -5.5
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"), -- 3.2 + -3.2 = 0
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000001000000000000000000000"), -- 2.6 + -0.1 = 2.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111110010011001100110011010000"), -- 3.5 + -3.7 = -0.2
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"00111110100110011001100110100000"), -- -3.1 + 3.4 = 0.3
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000100100000000000000000000"), -- -2.4 + -2.1 = -4.5
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111110110011001100110011001100"), -- 0.9 + -0.5 = 0.4
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000100011001100110011001101"), -- 1.2 + 3.2 = 4.4
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"10111111100011001100110011001101"), -- 1.4 + -2.5 = -1.1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000010011001100110011001101"), -- -0.7 + -2.5 = -3.2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000011001100110011001100111"), -- -0.3 + 3.9 = 3.6
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000100001100110011001100110"), -- 2.4 + 1.8 = 4.2
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000100011001100110011001101"), -- 1 + 3.4 = 4.4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000100101100110011001100110"), -- -3.8 + -0.9 = -4.7
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000001100110011001100110100"), -- -0.4 + -2.4 = -2.8
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000000001100110011001100111"), -- -0.8 + 2.9 = 2.1
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000000001000000000000000000000"), -- 3.3 + -0.8 = 2.5
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000001011001100110011001101"), -- 1 + -3.7 = -2.7
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000111000000000000000000000"), -- 3.9 + 3.1 = 7
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000101000000000000000000000"), -- 2.7 + 2.3 = 5
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000000011001100110011001101"), -- 1.3 + -3.5 = -2.2
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000000100110011001100110100"), -- 0.6 + 1.7 = 2.3
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111111111111111111111111111"), -- -2.6 + 0.6 = -2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111100000000000000000000000"), -- 0.2 + 0.8 = 1
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000100111001100110011001101"), -- 3.9 + 1 = 4.9
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111100011001100110011001100"), -- 2.7 + -3.8 = -1.1
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000010000000000000000000000"), -- 1 + 2 = 3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000000100110011001100110011"), -- 0.7 + -3 = -2.3
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000000001100110011001100110"), -- 0.5 + -2.6 = -2.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111111100110011001100110011010"), -- -1.2 + 2.4 = 1.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000010100110011001100110011"), -- -0.7 + -2.6 = -3.3
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"00111111010011001100110011001110"), -- 2.4 + -1.6 = 0.8
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000100101100110011001100110"), -- -1.3 + -3.4 = -4.7
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000001011001100110011001100"), -- 1.3 + 1.4 = 2.7
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111010011001100110011001101"), -- 0.8 + -1.6 = -0.8
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111000000000000000000000000"), -- -0.1 + -0.4 = -0.5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"10111111010011001100110011001101"), -- -0.7 + -0.1 = -0.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"10111110010011001100110011010000"), -- -2.8 + 2.6 = -0.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111101001100110011001100110"), -- -0.9 + -0.4 = -1.3
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111110100110011001100110011000"), -- 2.4 + -2.7 = -0.3
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000111100000000000000000000"), -- 3.9 + 3.6 = 7.5
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"10111110010011001100110011010000"), -- -1.6 + 1.4 = -0.2
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000010110011001100110011001"), -- 3.8 + -0.4 = 3.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111110010011001100110011010000"), -- -1.1 + 0.9 = -0.2
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000100001100110011001100110"), -- 1.9 + 2.3 = 4.2
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"10111111100000000000000000000000"), -- 1.7 + -2.7 = -1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"10111111011001100110011001100110"), -- 0 + -0.9 = -0.9
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111110011001100110011001101"), -- -1.4 + -0.2 = -1.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111110100110011001100110011000"), -- 3.3 + -3.6 = -0.3
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000110001100110011001100110"), -- 3.8 + 2.4 = 6.2
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111010011001100110011001100"), -- -0.1 + 0.9 = 0.8
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000000100110011001100110100"), -- -0.9 + 3.2 = 2.3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"), -- -2.5 + 2.5 = 0
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"10111111000110011001100110011000"), -- -3 + 2.4 = -0.6
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"10111101110011001100110011000000"), -- -2.6 + 2.5 = -0.0999999
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000100001100110011001100110"), -- -3.6 + -0.6 = -4.2
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"10111111001100110011001100110100"), -- -2.9 + 2.2 = -0.7
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111101001100110011001100110"), -- 1 + 0.3 = 1.3
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00111111110000000000000000000000"), -- 0 + 1.5 = 1.5
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000001001100110011001100110"), -- -3 + 0.4 = -2.6
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111111100011001100110011001101"), -- -1.6 + 2.7 = 1.1
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111110110011001100110011010000"), -- -3.2 + 2.8 = -0.4
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000100001100110011001100110"), -- -3.2 + -1 = -4.2
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"10111110010011001100110011010000"), -- -3.8 + 3.6 = -0.2
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111110011001100110011001100"), -- -2.2 + 3.8 = 1.6
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111111111100110011001100110100"), -- 2.2 + -0.3 = 1.9
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111010011001100110011001100"), -- -1.8 + 2.6 = 0.8
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100000110011001100110011"), -- 1 + 3.1 = 4.1
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000011001100110011001100110"), -- 2.6 + 1 = 3.6
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111111100110011001100110011"), -- 0.1 + 1.8 = 1.9
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000011011001100110011001101"), -- 0.5 + 3.2 = 3.7
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111000000000000000000000000"), -- 2.8 + -3.3 = -0.5
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"10111111110000000000000000000000"), -- -2 + 0.5 = -1.5
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111000000000000000000000000"), -- -0.5 + -0 = -0.5
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000101110011001100110011010"), -- -2.4 + -3.4 = -5.8
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000100000000000000000000000"), -- -3.5 + -0.5 = -4
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000001001100110011001100111"), -- -2.9 + 0.3 = -2.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000101101100110011001100110"), -- 2.7 + 3 = 5.7
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111011001100110011001101000"), -- 3.4 + -2.5 = 0.9
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000100001100110011001100110"), -- -3.3 + -0.9 = -4.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000100101100110011001100110"), -- 3.2 + 1.5 = 4.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"00111111000110011001100110011010"), -- 1.1 + -0.5 = 0.6
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"), -- 2.1 + -2.1 = 0
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"00111111110011001100110011001100"), -- 1.9 + -0.3 = 1.6
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"10111110010011001100110011010000"), -- 2.2 + -2.4 = -0.2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111111100110011001100110011010"), -- 2.4 + -1.2 = 1.2
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000010110011001100110011001"), -- -1.3 + -2.1 = -3.4
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"10111101110011001100110011010000"), -- -1.4 + 1.3 = -0.1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111101100110011001100110100"), -- 2.5 + -3.9 = -1.4
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000011011001100110011001100"), -- 1.8 + 1.9 = 3.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000011100110011001100110011"), -- 2.6 + 1.2 = 3.8
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111100011001100110011001110"), -- 2.8 + -3.9 = -1.1
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000100001100110011001100110"), -- -2.3 + -1.9 = -4.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + -0 = 0
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000010110011001100110011001"), -- -0.8 + -2.6 = -3.4
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000000110011001100110011010"), -- -0.3 + 2.7 = 2.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000001100110011001100110011"), -- 0.3 + -3.1 = -2.8
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000100000000000000000000000"), -- -0.8 + -3.2 = -4
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"10111111010011001100110011001100"), -- 1.1 + -1.9 = -0.8
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111101100110011001100110011"), -- -2.5 + 1.1 = -1.4
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000010011001100110011001100"), -- 2.6 + 0.6 = 3.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111000000000000000000000000"), -- -0.5 + 1 = 0.5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111100110011001100110011010"), -- -0.7 + -0.5 = -1.2
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"00111111111100110011001100110010"), -- 2.1 + -0.2 = 1.9
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111111100110011001100110100"), -- 1.7 + 0.2 = 1.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000000110011001100110011010"), -- 0 + -2.4 = -2.4
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010011001100110011001101"), -- 0.2 + -3.4 = -3.2
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111110010011001100110011010000"), -- -2 + 2.2 = 0.2
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"11000000000011001100110011001100"), -- -3.1 + 0.9 = -2.2
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111111001100110011001100110100"), -- -0.3 + -0.4 = -0.7
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000010011001100110011001101"), -- -2.5 + -0.7 = -3.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000001000000000000000000000"), -- -0.2 + 2.7 = 2.5
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"00111110010011001100110011001110"), -- -0.4 + 0.6 = 0.2
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111000110011001100110011010"), -- -0.6 + -0 = -0.6
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000001110011001100110011010"), -- -2.9 + -0 = -2.9
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000101000110011001100110011"), -- 2 + 3.1 = 5.1
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000011100110011001100110100"), -- -3.2 + -0.6 = -3.8
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000000000000000000000000000"), -- 1.7 + 0.3 = 2
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"10111111101100110011001100110011"), -- 0.2 + -1.6 = -1.4
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111111001100110011001100110"), -- -1 + -0.8 = -1.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000011001100110011001100110"), -- 0 + -3.6 = -3.6
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000011110011001100110011010"), -- 1.9 + 2 = 3.9
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000100011001100110011001101"), -- 0.7 + 3.7 = 4.4
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000011110011001100110011010"), -- 2.5 + 1.4 = 3.9
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111110011001100110011001100"), -- -2.8 + 1.2 = -1.6
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000011001100110011001100111"), -- -0.4 + -3.2 = -3.6
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"10111111011001100110011001100100"), -- 1.7 + -2.6 = -0.9
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000010000000000000000000000"), -- -3.4 + 0.4 = -3
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111000110011001100110011000"), -- -2.6 + 2 = -0.6
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000000100110011001100110011"), -- 2.3 + -0 = 2.3
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000001000000000000000000000"), -- 3.6 + -1.1 = 2.5
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111111110011001100110011001100"), -- 0.7 + -2.3 = -1.6
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000011001100110011001100110"), -- -3.1 + -0.5 = -3.6
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000000000001100110011001100110"), -- -0.8 + -1.3 = -2.1
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"00111111110000000000000000000000"), -- 2.8 + -1.3 = 1.5
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111110011001100110011001100"), -- -3.6 + 2 = -1.6
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"00111110110011001100110011010000"), -- -2.8 + 3.2 = 0.4
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000001100110011001100110100"), -- 1.2 + 1.6 = 2.8
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000011001100110011001100"), -- -3.6 + 1.4 = -2.2
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000101111001100110011001101"), -- -3.5 + -2.4 = -5.9
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000100000110011001100110011"), -- 0.3 + 3.8 = 4.1
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000001110011001100110011010"), -- 1.6 + 1.3 = 2.9
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000010110011001100110011010"), -- -1.8 + -1.6 = -3.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000110101100110011001100110"), -- 3 + 3.7 = 6.7
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000001001100110011001100110"), -- -3.8 + 1.2 = -2.6
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000000110011001100110011010"), -- -0.6 + -1.8 = -2.4
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"00111111111001100110011001100110"), -- 1.5 + 0.3 = 1.8
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000000100110011001100110100"), -- -1.1 + 3.4 = 2.3
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100100110011001100110011"), -- 1.1 + 3.5 = 4.6
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"00111110100110011001100110011000"), -- -2.9 + 3.2 = 0.3
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111111100110011001100110011000"), -- -2.4 + 3.6 = 1.2
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"10111111110110011001100110011010"), -- -3.2 + 1.5 = -1.7
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000011000000000000000000000"), -- 0.2 + 3.3 = 3.5
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111000000000000000000000000"), -- -2.8 + 3.3 = 0.5
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000000110011001100110011010"), -- -2.9 + 0.5 = -2.4
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000101100110011001100110011"), -- 1.9 + 3.7 = 5.6
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111111110011001100110011001110"), -- 2.1 + -3.7 = -1.6
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000000100110011001100110011"), -- 3 + -0.7 = 2.3
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000001011001100110011001100"), -- 1.4 + 1.3 = 2.7
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000000000000000000000000000"), -- 0.8 + 1.2 = 2
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111110100110011001100110011000"), -- -1.6 + 1.9 = 0.3
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000101100000000000000000000"), -- 3.7 + 1.8 = 5.5
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111111100110011001100110011001"), -- -3.1 + 1.9 = -1.2
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"00111111101001100110011001100111"), -- 0.1 + 1.2 = 1.3
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000100011001100110011001101"), -- -0.9 + -3.5 = -4.4
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101010011001100110011010"), -- -2.7 + -2.6 = -5.3
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000000001100110011001100111"), -- -1.8 + 3.9 = 2.1
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000000011011001100110011001101"), -- 3.4 + 0.3 = 3.7
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"10111111010011001100110011001110"), -- -1.7 + 0.9 = -0.8
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000101100110011001100110011"), -- 2.1 + 3.5 = 5.6
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000100011001100110011001101"), -- 0.9 + 3.5 = 4.4
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000111000000000000000000000"), -- 3.1 + 3.9 = 7
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000100000110011001100110011"), -- 2.3 + 1.8 = 4.1
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111100011001100110011001101"), -- -1.7 + 0.6 = -1.1
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111011001100110011001100110"), -- -0.4 + -0.5 = -0.9
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000100010011001100110011010"), -- 1.8 + 2.5 = 4.3
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000011000000000000000000000"), -- 3.5 + -0 = 3.5
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000010000000000000000000000"), -- 2.6 + 0.4 = 3
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111101001100110011001100111"), -- 1.6 + -2.9 = -1.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000000001100110011001100110"), -- 2.1 + -0 = 2.1
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000110011001100110011001101"), -- -2.5 + -3.9 = -6.4
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111010011001100110011001110"), -- -0.9 + 1.7 = 0.8
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"00111111110011001100110011001100"), -- -1.5 + 3.1 = 1.6
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111000110011001100110011100"), -- 2.8 + -3.4 = -0.6
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000010110011001100110011001"), -- -2.6 + -0.8 = -3.4
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000001110011001100110011010"), -- -0.4 + -2.5 = -2.9
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111111110110011001100110011010"), -- 3.8 + -2.1 = 1.7
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"00111111110011001100110011001100"), -- -0.5 + 2.1 = 1.6
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111010011001100110011001101"), -- 0.2 + -1 = -0.8
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000000001001100110011001100111"), -- 0.2 + 2.4 = 2.6
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000011011001100110011001101"), -- 3.7 + -0 = 3.7
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000001100110011001100110011"), -- -0.3 + 3.1 = 2.8
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111101110011001100110011000000"), -- -3.2 + 3.3 = 0.0999999
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111101100110011001100110100"), -- -0.8 + 2.2 = 1.4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"10111111110011001100110011001100"), -- -3.8 + 2.2 = -1.6
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000001000000000000000000000"), -- 3.6 + -1.1 = 2.5
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000100000110011001100110011"), -- -3 + -1.1 = -4.1
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"00111111100011001100110011001100"), -- 3.8 + -2.7 = 1.1
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000101100110011001100110100"), -- 2.7 + 2.9 = 5.6
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000100011001100110011001101"), -- -1.5 + -2.9 = -4.4
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"00111111100110011001100110011010"), -- 3.7 + -2.5 = 1.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111111000110011001100110011010"), -- -0.5 + 1.1 = 0.6
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000010011001100110011001101"), -- 2.8 + 0.4 = 3.2
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111011001100110011001100110"), -- 1 + -0.1 = 0.9
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000111000110011001100110100"), -- -3.9 + -3.2 = -7.1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111110000000000000000000000"), -- 0.6 + 0.9 = 1.5
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000001000000000000000000000"), -- -1 + 3.5 = 2.5
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000100110011001100110011010"), -- -2.9 + -1.9 = -4.8
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000101101100110011001100110"), -- 1.8 + 3.9 = 5.7
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111110010011001100110011001100"), -- 0.6 + -0.8 = -0.2
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000110010011001100110011010"), -- -3.7 + -2.6 = -6.3
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111100000000000000000000000"), -- 0.8 + 0.2 = 1
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000001100110011001100110011"), -- -1.8 + -1 = -2.8
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111101110011001100110011010000"), -- 1.1 + -1.2 = -0.1
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000000000000000000000000000"), -- -3.4 + 1.4 = -2
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000010011001100110011001101"), -- 0.4 + 2.8 = 3.2
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000101100110011001100110100"), -- -3.9 + -1.7 = -5.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000000100110011001100110011"), -- -1.3 + -1 = -2.3
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000010000000000000000000000"), -- -2.5 + -0.5 = -3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111111111100110011001100110100"), -- -0.5 + 2.4 = 1.9
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000100001100110011001100110"), -- -0.5 + -3.7 = -4.2
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000101001100110011001100110"), -- -1.7 + -3.5 = -5.2
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000100011001100110011001101"), -- 1 + 3.4 = 4.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000100100000000000000000000"), -- -1.1 + -3.4 = -4.5
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111110110011001100110011010000"), -- 2.2 + -1.8 = 0.4
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111111101001100110011001100110"), -- 0.7 + -2 = -1.3
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000011000000000000000000000"), -- 2.5 + 1 = 3.5
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"00111110110011001100110011001100"), -- 1.6 + -1.2 = 0.4
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111111100110011001100110011010"), -- -1.9 + 0.7 = -1.2
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111101001100110011001100110"), -- 2.3 + -3.6 = -1.3
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111100000000000000000000001"), -- 2.9 + -1.9 = 1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"00111111100110011001100110011010"), -- -0.8 + 2 = 1.2
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111111001100110011001100110010"), -- 1.8 + -1.1 = 0.7
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111000000000000000000000000"), -- -1.3 + 1.8 = 0.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010000000000000000000000"), -- 0.4 + -3.4 = -3
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000100100000000000000000000"), -- 2 + 2.5 = 4.5
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111101100110011001100110100"), -- -0.3 + 1.7 = 1.4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000010001100110011001100111"), -- 2.7 + 0.4 = 3.1
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000100101100110011001100110"), -- -3.6 + -1.1 = -4.7
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"10111111110110011001100110011010"), -- -3 + 1.3 = -1.7
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111111000000000000000000000000"), -- -2.2 + 2.7 = 0.5
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111110011001100110011001100"), -- 1.2 + -2.8 = -1.6
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111101110011001100110011000000"), -- -3.4 + 3.5 = 0.0999999
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111110011001100110011001101"), -- -1.4 + -0.2 = -1.6
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"10111111111001100110011001100110"), -- 0.7 + -2.5 = -1.8
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"10111111110000000000000000000000"), -- -3.7 + 2.2 = -1.5
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"00111111110011001100110011001110"), -- -2.3 + 3.9 = 1.6
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"10111111110000000000000000000000"), -- -2.2 + 0.7 = -1.5
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000010110011001100110011010"), -- 3.7 + -0.3 = 3.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101010011001100110011010"), -- -3.7 + -1.6 = -5.3
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00111111101111111111111111111111"), -- 2.1 + -0.6 = 1.5
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111111010011001100110011001101"), -- 1.5 + -0.7 = 0.8
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000100101100110011001100110"), -- 2.2 + 2.5 = 4.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000011001100110011001100110"), -- 2.6 + 1 = 3.6
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000001000000000000000000000"), -- 3.6 + -1.1 = 2.5
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000000011001100110011001100"), -- 1.3 + 0.9 = 2.2
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"00111111110000000000000000000000"), -- 3.7 + -2.2 = 1.5
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111110100110011001100110011000"), -- 2.7 + -2.4 = 0.3
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000011000000000000000000000"), -- -1.3 + -2.2 = -3.5
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000010110011001100110011010"), -- 0 + -3.4 = -3.4
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111100110011001100110011010"), -- 0.2 + 1 = 1.2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111110110011001100110011001000"), -- 2.4 + -2.8 = -0.4
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000011110011001100110011010"), -- 0.4 + 3.5 = 3.9
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000010110011001100110011010"), -- -2.3 + -1.1 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111010011001100110011001101"), -- 0 + -0.8 = -0.8
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000010100110011001100110011"), -- 3.3 + -0 = 3.3
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000101001100110011001100110"), -- 1.9 + 3.3 = 5.2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111101110011001100110011010000"), -- -1.2 + 1.1 = -0.1
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000111001100110011001100110"), -- 3.9 + 3.3 = 7.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111110000000000000000000000"), -- -0.9 + -0.6 = -1.5
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000110100110011001100110100"), -- -2.9 + -3.7 = -6.6
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111000110011001100110011000"), -- -2.2 + 2.8 = 0.6
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111000110011001100110011010"), -- -1.1 + 1.7 = 0.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000100111001100110011001101"), -- -2 + -2.9 = -4.9
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111111001100110011001100110"), -- 1.3 + 0.5 = 1.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000011001100110011001100111"), -- 3.9 + -0.3 = 3.6
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000110000000000000000000000"), -- -2.4 + -3.6 = -6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"00111110110011001100110011001101"), -- 0.8 + -0.4 = 0.4
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111110100110011001100110011000"), -- 2.8 + -3.1 = -0.3
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"10111111111111111111111111111111"), -- -2.1 + 0.1 = -2
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000101100110011001100110011"), -- -1.8 + -3.8 = -5.6
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000011001100110011001100110"), -- -1.9 + -1.7 = -3.6
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"10111111000110011001100110011000"), -- -3 + 2.4 = -0.6
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000100000110011001100110011"), -- -0.4 + -3.7 = -4.1
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000100000000000000000000000"), -- 2.6 + 1.4 = 4
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111100110011001100110011010"), -- -0.1 + -1.1 = -1.2
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110100110011001100110100"), -- -3.7 + -2.9 = -6.6
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000000011001100110011001100"), -- 1.1 + -3.3 = -2.2
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000000110011001100110011010"), -- -2.9 + 0.5 = -2.4
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000010100110011001100110011"), -- -1.5 + -1.8 = -3.3
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111110110011001100110011001"), -- 1.8 + -0.1 = 1.7
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000100000000000000000000000"), -- 3.1 + 0.9 = 4
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000010100110011001100110011"), -- 1 + 2.3 = 3.3
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000000100110011001100110011"), -- 2.2 + 0.1 = 2.3
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000011001100110011001100110"), -- 2 + 1.6 = 3.6
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000101010011001100110011010"), -- 3.4 + 1.9 = 5.3
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111000110011001100110011010"), -- 2.5 + -1.9 = 0.6
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000000110011001100110011010"), -- 2.5 + -0.1 = 2.4
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000001000000000000000000000"), -- -0.5 + 3 = 2.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"00111111000110011001100110011010"), -- 2.5 + -1.9 = 0.6
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000110100000000000000000000"), -- -3.8 + -2.7 = -6.5
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"00111111100000000000000000000000"), -- -0.7 + 1.7 = 1
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"10111101110011001100110011000000"), -- -3.3 + 3.2 = -0.0999999
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111000000000000000000000000"), -- -3.3 + 3.8 = 0.5
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000110101100110011001100110"), -- -3.2 + -3.5 = -6.7
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000011000000000000000000000"), -- 2.5 + 1 = 3.5
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"10111111100011001100110011001100"), -- -3.3 + 2.2 = -1.1
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"10111111101001100110011001100110"), -- 1 + -2.3 = -1.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101000000000000000000000"), -- 2.8 + 2.2 = 5
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"00111111100011001100110011001101"), -- -0.9 + 2 = 1.1
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000011100110011001100110011"), -- -0.5 + -3.3 = -3.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"00111111110000000000000000000000"), -- 3.7 + -2.2 = 1.5
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000010100110011001100110011"), -- 3.7 + -0.4 = 3.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"10111111100000000000000000000000"), -- -1 + -0 = -1
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110101100110011001100110"), -- -3.8 + -2.9 = -6.7

	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000000111111111111111111111"), -- -1.7 + 4.2 = 2.5
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000110011001100110011001100"), -- -5.2 + -1.2 = -6.4
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001011011100110011001100110"), -- -5.9 + -9 = -14.9
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000000101001100110011001100111"), -- -0.2 + 5.4 = 5.2
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"01000000100101100110011001100110"), -- -1.3 + 6 = 4.7
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"10111111000000000000000000000000"), -- -9.4 + 8.9 = -0.5
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000100000000000000000000", b"01000001011000000000000000000000"), -- 5 + 9 = 14
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000000110100110011001100110100"), -- 1.7 + 4.9 = 6.6
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000001000101100110011001100110"), -- -6 + -3.4 = -9.4
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"10111111101001100110011001100110"), -- -1.9 + 0.6 = -1.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000001111111111111111111111"), -- -1.2 + 4.2 = 3
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000001001110000000000000000000"), -- -5 + -6.5 = -11.5
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000100110011001100110011010"), -- 6.5 + -1.7 = 4.8
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000001000011001100110011001101"), -- 7.6 + 1.2 = 8.8
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000001100000100110011001100110"), -- 9.8 + 6.5 = 16.3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000000000000000000000000000"), -- 0.7 + 1.3 = 2
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"11000001010101100110011001100110"), -- -6.4 + -7 = -13.4
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000000100101100110011001100110"), -- 4.5 + -9.2 = -4.7
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"00111111110000000000000000000000"), -- 9.2 + -7.7 = 1.5
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000000110101100110011001100111"), -- -0.4 + -6.3 = -6.7
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"00111111101100110011001100110100"), -- -4.5 + 5.9 = 1.4
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000001010101001100110011001100"), -- -9.9 + -3.4 = -13.3
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000100111001100110011001100"), -- 3.1 + 1.8 = 4.9
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"00111111000110011001100110011000"), -- 5 + -4.4 = 0.6
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111100110011001100110011010"), -- 2.1 + -3.3 = -1.2
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"01000000100000110011001100110011"), -- -1.9 + 6 = 4.1
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"01000000101110011001100110011001"), -- 9.2 + -3.4 = 5.8
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000000001000000000000000000010"), -- 7.1 + -9.6 = -2.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"11000000111110011001100110011010"), -- -0 + -7.8 = -7.8
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000000111110011001100110011001"), -- 1.1 + 6.7 = 7.8
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000001000110000000000000000000"), -- -4.1 + -5.4 = -9.5
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"10111111000110011001100110011000"), -- -7 + 6.4 = -0.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00111110110011001100110011010000"), -- -2 + 2.4 = 0.4
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"01000000111110011001100110011010"), -- 1.9 + 5.9 = 7.8
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"10111110110011001100110011000000"), -- 9.5 + -9.9 = -0.4
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000010000000000000000000000"), -- 1.9 + 1.1 = 3
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"11000000101101100110011001100110"), -- -9.5 + 3.8 = -5.7
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001000000000000000000000"), -- 2.7 + -0.2 = 2.5
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000000100000110011001100110011"), -- 2.1 + -6.2 = -4.1
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100101100110011001100110", b"00111111100011001100110011010000"), -- 5.8 + -4.7 = 1.1
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000001000100110011001100110011"), -- -6.7 + -2.5 = -9.2
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"00111111101100110011001100110000"), -- -5.3 + 6.7 = 1.4
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111000110011001100110011100"), -- 2.8 + -3.4 = -0.6
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000001000011001100110011001101"), -- -5.6 + -3.2 = -8.8
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"10111111110011001100110011010000"), -- 4.7 + -6.3 = -1.6
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000000101100000000000000000000"), -- 6.4 + -0.9 = 5.5
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101100000000000000000000", b"01000001011010000000000000000000"), -- 9 + 5.5 = 14.5
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001001010000000000000000000"), -- 4.4 + 6.1 = 10.5
	(b"11000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000001010100000000000000000000"), -- -8.8 + -4.2 = -13
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"01000000101000000000000000000000"), -- 8.3 + -3.3 = 5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000000101100110011001100110011"), -- -0 + -5.6 = -5.6
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"01000000110000000000000000000000"), -- 8 + -2 = 6
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001100010001100110011001101"), -- -7.6 + -9.5 = -17.1
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001001111001100110011001100"), -- -2.9 + -8.9 = -11.8
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"01000001010010011001100110011010"), -- 5.1 + 7.5 = 12.6
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"10111111111001100110011001100110"), -- -5 + 3.2 = -1.8
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"00111111010011001100110011000000"), -- -8.6 + 9.4 = 0.799999
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"01000000011000000000000000000000"), -- -4 + 7.5 = 3.5
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000001001101100110011001100110"), -- 8.5 + 2.9 = 11.4
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000001011001001100110011001101"), -- 9 + 5.3 = 14.3
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"10111111100011001100110011001100"), -- -3.1 + 2 = -1.1
	(b"01000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000001000011001100110011001101"), -- 6.6 + 2.2 = 8.8
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"11000000110111001100110011001101"), -- -8 + 1.1 = -6.9
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000111010011001100110011010"), -- 5.4 + 1.9 = 7.3
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000001011100110011001100110100"), -- 7.9 + 7.3 = 15.2
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000111001100110011001100111"), -- 7.9 + -0.7 = 7.2
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000101011001100110011001101"), -- 3.9 + 1.5 = 5.4
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000001000000000000000000000"), -- -2.1 + -0.4 = -2.5
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"11000001011000011001100110011010"), -- -7.2 + -6.9 = -14.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000000100100110011001100110100"), -- -1.2 + 5.8 = 4.6
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000001000010110011001100110011"), -- 8.3 + 0.4 = 8.7
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"01000000000011001100110011001100"), -- 6.1 + -3.9 = 2.2
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000001001010110011001100110011"), -- -7.6 + -3.1 = -10.7
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"01000000110001100110011001100111"), -- 7.8 + -1.6 = 6.2
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000000111100000000000000000000"), -- 3.4 + 4.1 = 7.5
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000000011001100110011001100111"), -- -4.9 + 1.3 = -3.6
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001010110000000000000000000"), -- 4 + 9.5 = 13.5
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000000111101100110011001100110"), -- -1.7 + -6 = -7.7
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"01000000100010011001100110011010"), -- -0.2 + 4.5 = 4.3
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"11000000110101100110011001100111"), -- -8.6 + 1.9 = -6.7
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000001001111001100110011001100"), -- -9.4 + -2.4 = -11.8
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000001100011001100110011001100"), -- 8.7 + 8.9 = 17.6
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000000100101100110011001100110"), -- 3.7 + -8.4 = -4.7
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000001010101100110011001100110"), -- 4.7 + 8.7 = 13.4
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000001000100011001100110011010"), -- 7 + 2.1 = 9.1
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000001000100011001100110011010"), -- -8.3 + -0.8 = -9.1
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000101000000000000000000000"), -- -2.2 + 7.2 = 5
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000001011000110011001100110011"), -- 8.5 + 5.7 = 14.2
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"01000000110000110011001100110011"), -- 2.1 + 4 = 6.1
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001100100110011001100110011"), -- -9 + -9.4 = -18.4
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000001000011100110011001100110"), -- 6.9 + 2 = 8.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"), -- 0 + 0 = 0
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- 0 + -2.8 = -2.8
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"10111110100110011001100110011000"), -- -4 + 3.7 = -0.3
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"00111111101100110011001100110100"), -- 9.3 + -7.9 = 1.4
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000001010000000000000000000000"), -- -7 + -5 = -12
	(b"11000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001011000000000000000000000"), -- -8.8 + -5.2 = -14
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000000100100000000000000000000"), -- 1.4 + -5.9 = -4.5
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001000000110011001100110011"), -- -0.2 + -8 = -8.2
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001010010110011001100110011"), -- -3 + -9.7 = -12.7
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000000101100110011001100110100"), -- 0.3 + 5.3 = 5.6
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"11000000100001100110011001100110"), -- -7.4 + 3.2 = -4.2
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000001010000000000000000000000"), -- 9.3 + 2.7 = 12
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000010001100110011001100110"), -- -0.6 + 3.7 = 3.1
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000001000111001100110011001101"), -- 1.9 + 7.9 = 9.8
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000000001110011001100110011010"), -- 6.4 + -9.3 = -2.9
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001011010000000000000000000"), -- -5.8 + -8.7 = -14.5
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000110011001100110011001101"), -- -3.9 + -2.5 = -6.4
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001010010000000000000000000"), -- -7.6 + -4.9 = -12.5
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000001010010110011001100110011"), -- 4.2 + 8.5 = 12.7
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"10111111111100110011001100110100"), -- -6.6 + 4.7 = -1.9
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000001010000000000000000000000"), -- -9.3 + -2.7 = -12
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000101011001100110011001101"), -- -0.6 + -4.8 = -5.4
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"11000001011011001100110011001101"), -- -5.7 + -9.1 = -14.8
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"00111111000110011001100110011000"), -- -7.9 + 8.5 = 0.6
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000100100000000000000000000"), -- -3.3 + -1.2 = -4.5
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001001000000000000000000000"), -- -1.8 + -8.2 = -10
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000000100101100110011001100111"), -- -2.1 + 6.8 = 4.7
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000000100100000000000000000000"), -- -3.1 + 7.6 = 4.5
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000111010011001100110011010"), -- -6.4 + -0.9 = -7.3
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000110001100110011001100110"), -- 7.2 + -1 = 6.2
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111111011001100110011001100110"), -- 0.4 + 0.5 = 0.9
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000001001011001100110011001100"), -- -7.2 + -3.6 = -10.8
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"01000001100100011001100110011010"), -- 9.9 + 8.3 = 18.2
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000000000100110011001100110011"), -- 3.7 + -6 = -2.3
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000000000000000000000000000"), -- 0.5 + 1.5 = 2
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001001111100110011001100110"), -- -3 + -8.9 = -11.9
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001011100011001100110011010"), -- -5.4 + -9.7 = -15.1
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000001000011001100110011001100"), -- 4.7 + 4.1 = 8.8
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001011100110011001100110011"), -- -8.9 + -6.3 = -15.2
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000000000001100110011001100110"), -- 2.9 + -5 = -2.1
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"01000000001110011001100110011010"), -- 5.4 + -2.5 = 2.9
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000001001010000000000000000000"), -- -4.6 + -5.9 = -10.5
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001011100110011001100110011"), -- -7.7 + -7.5 = -15.2
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001000011001100110011001100"), -- -3.6 + -5.2 = -8.8
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000001001100110011001100111"), -- 4.3 + -1.7 = 2.6
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000001001011100110011001100110"), -- 7 + 3.9 = 10.9
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000110010011001100110011001"), -- -7.7 + 1.4 = -6.3
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"11000000100000000000000000000000"), -- -7.4 + 3.4 = -4
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000001001101001100110011001100"), -- 7.2 + 4.1 = 11.3
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000110010011001100110011001"), -- 6.7 + -0.4 = 6.3
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000100110011001100110011010"), -- -5 + 0.2 = -4.8
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000001000010000000000000000000"), -- -0.9 + 9.4 = 8.5
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"10111111110000000000000000000000"), -- 4.1 + -5.6 = -1.5
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000001011110110011001100110100"), -- 8.1 + 7.6 = 15.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000010000000000000000000000"), -- 2.6 + 0.4 = 3
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001010110110011001100110011"), -- 7.6 + 6.1 = 13.7
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111010011001100110011001100"), -- -2.7 + 3.5 = 0.8
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000000110000000000000000000000"), -- 0.8 + 5.2 = 6
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000100010011001100110011010"), -- 6 + -1.7 = 4.3
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000001011111100110011001100110"), -- 7.1 + 8.8 = 15.9
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"00111111100110011001100110011001"), -- 2.1 + -0.9 = 1.2
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000001000101001100110011001101"), -- -8.2 + -1.1 = -9.3
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000001100011011001100110011010"), -- 9.3 + 8.4 = 17.7
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000000010100110011001100110010"), -- 6.4 + -9.7 = -3.3
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000001000010011001100110011010"), -- 1.2 + 7.4 = 8.6
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"11000001010100011001100110011010"), -- -6.1 + -7 = -13.1
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001001010110011001100110100"), -- -5.8 + -4.9 = -10.7
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"11000000010000000000000000000000"), -- -9.7 + 6.7 = -3
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000001001110110011001100110011"), -- 4 + 7.7 = 11.7
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"10111111010011001100110011010000"), -- 5 + -5.8 = -0.8
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000111111001100110011001100"), -- 9.4 + -1.5 = 7.9
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"11000001100100000000000000000000"), -- -8.9 + -9.1 = -18
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11000000101110011001100110011010"), -- -5.8 + 0 = -5.8
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000100100000000000000000000"), -- -0.7 + -3.8 = -4.5
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"01000000111010011001100110011001"), -- 9.9 + -2.6 = 7.3
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000001010100011001100110011010"), -- -9.5 + -3.6 = -13.1
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"01000001001011100110011001100110"), -- 5 + 5.9 = 10.9
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000001000100110011001100110100"), -- 4.3 + 4.9 = 9.2
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000100000000000000000000000"), -- 2.6 + 1.4 = 4
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001100010100110011001100110"), -- -8.6 + -8.7 = -17.3
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000000101111001100110011001100"), -- -4 + 9.9 = 5.9
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000100111001100110011001101"), -- -5.9 + 1 = -4.9
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001000011001100110011001101"), -- 1.8 + 7 = 8.8
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000001011100110011001100110011"), -- 9.4 + 5.8 = 15.2
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111111101100110011001100110011"), -- 0 + -1.4 = -1.4
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000000111100110011001100110011"), -- -1.9 + 9.5 = 7.6
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001001010110011001100110011"), -- 6.5 + 4.2 = 10.7
	(b"11000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"00111111100110011001100110100000"), -- -8.4 + 9.6 = 1.2
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001010101100110011001100111"), -- 3.8 + 9.6 = 13.4
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000000110001100110011001100111"), -- -0.8 + -5.4 = -6.2
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000000101101100110011001100111"), -- 1.6 + -7.3 = -5.7
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"01000000010000000000000000000000"), -- 7.3 + -4.3 = 3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"01000000111010011001100110011010"), -- 0.9 + 6.4 = 7.3
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"11000000101000000000000000000000"), -- -8 + 3 = -5
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000001000010110011001100110011"), -- -4.5 + -4.2 = -8.7
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"00111111011001100110011001100111"), -- 0.1 + 0.8 = 0.9
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"10111111000110011001100110100000"), -- -6.8 + 6.2 = -0.6
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11000000001011001100110011001101"), -- -2.7 + 0 = -2.7
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000010011001100110011001100"), -- -1 + 4.2 = 3.2
	(b"01000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"01000000110010011001100110011010"), -- 8.6 + -2.3 = 6.3
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001001001100110011001100110"), -- -4.7 + -5.7 = -10.4
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000000010001100110011001100110"), -- 4.9 + -8 = -3.1
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"11000000100011001100110011001100"), -- -7.1 + 2.7 = -4.4
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000100011001100110011001101"), -- 4.6 + -0.2 = 4.4
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000011110011001100110011010"), -- 4 + -0.1 = 3.9
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000101111001100110011001101"), -- -6.1 + 0.2 = -5.9
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"10111111000110011001100110011010"), -- 0.5 + -1.1 = -0.6
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"01000000011000000000000000000000"), -- 6.9 + -3.4 = 3.5
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000001000111001100110011001101"), -- 7.1 + 2.7 = 9.8
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"01000000101000000000000000000000"), -- 9.2 + -4.2 = 5
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000111110011001100110011010"), -- -4.6 + -3.2 = -7.8
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000010100110011001100110100"), -- 1.1 + 2.2 = 3.3
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000110010011001100110011010"), -- 3 + 3.3 = 6.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001000010011001100110011010"), -- -1 + 9.6 = 8.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000000101000000000000000000000"), -- 3.5 + -8.5 = -5
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100010011001100110011010", b"11000000000011001100110011001100"), -- -6.5 + 4.3 = -2.2
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"00111110100110011001100110100000"), -- -5.7 + 6 = 0.3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"10111111111001100110011001101000"), -- 2.6 + -4.4 = -1.8
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000001000010110011001100110011"), -- 8 + 0.7 = 8.7
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"00111110010011001100110011000000"), -- -9.3 + 9.5 = 0.2
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000100110011001100110011010"), -- -2.8 + -2 = -4.8
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000001000011100110011001100110"), -- -2.2 + -6.7 = -8.9
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001000110110011001100110011"), -- -1.5 + -8.2 = -9.7
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"11000000110011001100110011001101"), -- 0.5 + -6.9 = -6.4
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000011001100110011001100110"), -- 3.8 + -0.2 = 3.6
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000001001100011001100110011010"), -- 8.3 + 2.8 = 11.1
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"10111111000110011001100110010000"), -- -9.9 + 9.3 = -0.599999
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000000100111001100110011001101"), -- 4.4 + -9.3 = -4.9
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111111100110011001100110100"), -- 4.3 + -2.4 = 1.9
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"11000000101110011001100110011001"), -- -9.2 + 3.4 = -5.8
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000000110000000000000000000000"), -- -1.1 + -4.9 = -6
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"), -- 4 + -4 = 0
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000110010011001100110011010"), -- 4.8 + 1.5 = 6.3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000000111001100110011001100110"), -- 0.7 + 6.5 = 7.2
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000111011001100110011001101"), -- 5.8 + 1.6 = 7.4
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"00111111011111111111111111111111"), -- -0.8 + 1.8 = 1
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000000100011001100110011001100"), -- -0.8 + 5.2 = 4.4
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000100100000000000000000000"), -- 4.5 + -0 = 4.5
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000000111100000000000000000000"), -- -1.3 + -6.2 = -7.5
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"11000001001000110011001100110011"), -- -6.2 + -4 = -10.2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000000100101100110011001100111"), -- 0.7 + -5.4 = -4.7
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001001001100110011001100110"), -- -5.9 + -4.5 = -10.4
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000001100110001100110011001101"), -- 9.3 + 9.8 = 19.1
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000000001000000000000000000000"), -- 7.2 + -9.7 = -2.5
	(b"01000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"), -- 8.2 + -8.2 = 0
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"10111110010011001100110011001000"), -- 1.2 + -1.4 = -0.2
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111100000000000000000000000"), -- 0.8 + 0.2 = 1
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000001000000000000000000000000"), -- 4.4 + 3.6 = 8
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001001000011001100110011010"), -- -0.6 + -9.5 = -10.1
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"10111111000110011001100110100000"), -- -9 + 8.4 = -0.6
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000111010011001100110011010"), -- -7.3 + -0 = -7.3
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"10111111100110011001100110011001"), -- 1.9 + -3.1 = -1.2
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"11000000001100110011001100110011"), -- -5.5 + 2.7 = -2.8
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"11000001000111001100110011001100"), -- -4.7 + -5.1 = -9.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000000011110011001100110011010"), -- 3.9 + 0 = 3.9
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000001000110011001100110011010"), -- 7.4 + 2.2 = 9.6
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"01000000100000110011001100110100"), -- 7.8 + -3.7 = 4.1
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000010000000000000000000000"), -- -3.7 + 0.7 = -3
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001100000110011001100110011"), -- -8.2 + -8.2 = -16.4
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001000110000000000000000000"), -- 2.5 + 7 = 9.5
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000000001110011001100110011010"), -- 6.1 + -9 = -2.9
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000001100001001100110011001101"), -- 7.3 + 9.3 = 16.6
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000000001100110011001100110010"), -- 6.4 + -9.2 = -2.8
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000001000100000000000000000000"), -- 3.2 + 5.8 = 9
	(b"01000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"01000000000001100110011001100110"), -- 8.2 + -6.1 = 2.1
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111111011001100110011001100111"), -- -1.1 + 0.2 = -0.9
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"00111111101100110011001100110100"), -- 6.8 + -5.4 = 1.4
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000101000110011001100110011"), -- -2.3 + -2.8 = -5.1
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000001010010110011001100110100"), -- -6.8 + -5.9 = -12.7
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000100000000000000000000000"), -- -2.9 + -1.1 = -4
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"10111111111001100110011001101000"), -- 3.6 + -5.4 = -1.8
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"00111111001100110011001100110000"), -- 9.3 + -8.6 = 0.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000001000101001100110011001100"), -- 2.6 + 6.7 = 9.3
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000001011100110011001100110011"), -- 7.6 + 7.6 = 15.2
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"10111111011001100110011001100000"), -- 9 + -9.9 = -0.9
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000001010000110011001100110011"), -- 4.6 + 7.6 = 12.2
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"01000000101011001100110011001101"), -- -2.1 + 7.5 = 5.4
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"11000000100101100110011001100110"), -- -6.5 + 1.8 = -4.7
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000000000000000000000000000000"), -- -5.7 + 7.7 = 2
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"11000000001000000000000000000000"), -- -3.6 + 1.1 = -2.5
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000001000100000000000000000000"), -- -2.8 + -6.2 = -9
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000000010110011001100110011010"), -- -2 + 5.4 = 3.4
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000111010011001100110011001"), -- -7.6 + 0.3 = -7.3
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"10111111110011001100110011001100"), -- -7 + 5.4 = -1.6
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000001010111100110011001100110"), -- -9.5 + -4.4 = -13.9
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000000111101100110011001100110"), -- -1.8 + 9.5 = 7.7
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000001011001001100110011001100"), -- -5.1 + -9.2 = -14.3
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000001000100110011001100110011"), -- 9.7 + -0.5 = 9.2
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000001100011100110011001100110"), -- -8.5 + -9.3 = -17.8
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"00111111101001100110011001100100"), -- 4.7 + -3.4 = 1.3
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001000000000000000000000000"), -- -0.4 + -7.6 = -8
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"01000000001011001100110011001100"), -- 4.1 + -1.4 = 2.7
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000001010000110011001100110100"), -- -3.4 + -8.8 = -12.2
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000010100110011001100110011"), -- -3.5 + 0.2 = -3.3
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000001010011001100110011001100"), -- 6.1 + 6.7 = 12.8
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000001010110110011001100110100"), -- -5.1 + -8.6 = -13.7
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000011110011001100110011010"), -- -3 + -0.9 = -3.9
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000001100110001100110011001100"), -- -9.2 + -9.9 = -19.1
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"01000001001101100110011001100110"), -- 6.9 + 4.5 = 11.4
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000001011101100110011001100110"), -- 9.2 + 6.2 = 15.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111011001100110011001101", b"11000000111011001100110011001101"), -- 0 + -7.4 = -7.4
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000001001100110011001100110011"), -- 7.9 + 3.3 = 11.2
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000001000010011001100110011001"), -- -8.7 + 0.1 = -8.6
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000100101100110011001100110"), -- -2.5 + -2.2 = -4.7
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000000100011001100110011001100"), -- -2.3 + 6.7 = 4.4
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000110001100110011001100111"), -- 5.4 + 0.8 = 6.2
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000001100011110011001100110100"), -- 8.1 + 9.8 = 17.9
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"00111111011001100110011001100000"), -- 9.9 + -9 = 0.9
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"10111111101001100110011001101000"), -- 5 + -6.3 = -1.3
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001001110110011001100110011"), -- -7.2 + -4.5 = -11.7
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000000110111001100110011001110"), -- -2.7 + 9.6 = 6.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000000110001100110011001100110"), -- -0.9 + 7.1 = 6.2
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000010110011001100110011001"), -- 0.1 + 3.3 = 3.4
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000001100110100110011001100110"), -- -9.7 + -9.6 = -19.3
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000001000101001100110011001101"), -- 0.5 + -9.8 = -9.3
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"10111110100110011001100110100000"), -- -6.8 + 6.5 = -0.3
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000001000001001100110011001101"), -- -6 + -2.3 = -8.3
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"10111111110011001100110011001100"), -- -5.1 + 3.5 = -1.6
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000100010011001100110011010"), -- 0.4 + 3.9 = 4.3
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000110100110011001100110011"), -- 6.4 + 0.2 = 6.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"00111111001100110011001100110011"), -- 1.5 + -0.8 = 0.7
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000000011001100110011001100111"), -- 1.8 + -5.4 = -3.6
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000000011110011001100110011010"), -- -4.9 + 8.8 = 3.9
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000001001101001100110011001100"), -- 5.6 + 5.7 = 11.3
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000000000011001100110011001110"), -- -6.9 + 9.1 = 2.2
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000000010001100110011001100111"), -- -2.7 + 5.8 = 3.1
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"01000000110011001100110011001100"), -- 8.7 + -2.3 = 6.4
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"00111111110110011001100110011000"), -- 6.5 + -4.8 = 1.7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"11000000010100110011001100110011"), -- 3.7 + -7 = -3.3
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"00111110010011001100110011000000"), -- 8.7 + -8.5 = 0.2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"10111111101001100110011001100110"), -- 2.4 + -3.7 = -1.3
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"00111101110011001100110011000000"), -- 4.9 + -4.8 = 0.0999999
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000000101001100110011001100111"), -- 2.1 + -7.3 = -5.2
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000001000111100110011001100110"), -- 4.5 + 5.4 = 9.9
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000001010011100110011001100110"), -- -5.2 + -7.7 = -12.9
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000001000010011001100110011010"), -- -4.5 + -4.1 = -8.6
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"00111111111001100110011001101000"), -- -4 + 5.8 = 1.8
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000110100000000000000000000"), -- -4.7 + -1.8 = -6.5
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000001001011100110011001100111"), -- -9.1 + -1.8 = -10.9
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000101100110011001100110011"), -- -6.6 + 1 = -5.6
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000101011001100110011001101"), -- -4.3 + -1.1 = -5.4
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000101001100110011001100110"), -- 1.5 + 3.7 = 5.2
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001001011100110011001100110"), -- -2.7 + -8.2 = -10.9
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000000000110011001100110011000"), -- 5.3 + -7.7 = -2.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000011110011001100110011001"), -- -3.3 + 7.2 = 3.9
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000001010000011001100110011010"), -- 9.2 + 2.9 = 12.1
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000001000011100110011001100110"), -- -7.9 + -1 = -8.9
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"10111111010011001100110011010000"), -- -4.3 + 3.5 = -0.8
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111111000000000000000000000000"), -- 2.3 + -1.8 = 0.5
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000000000000000000000000000"), -- -0.2 + 2.2 = 2
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"10111111100000000000000000000000"), -- -9.9 + 8.9 = -1
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000001011011001100110011001101"), -- 8.5 + 6.3 = 14.8
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"10111111100011001100110011001100"), -- 5.4 + -6.5 = -1.1
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100101100110011001100110", b"01000000000000000000000000000000"), -- 6.7 + -4.7 = 2
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"01000000110011001100110011001101"), -- 1.4 + 5 = 6.4
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000111000110011001100110011"), -- 5 + 2.1 = 7.1
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000001010101001100110011001101"), -- 9.6 + 3.7 = 13.3
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001000101100110011001100110"), -- -4.1 + -5.3 = -9.4
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"11000000101100000000000000000000"), -- -9.2 + 3.7 = -5.5
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000001100000100110011001100110"), -- -9.6 + -6.7 = -16.3
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"00111111010011001100110011010000"), -- 4.9 + -4.1 = 0.8
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000100000110011001100110011"), -- -2 + -2.1 = -4.1
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001010110011001100110011010"), -- 4 + 9.6 = 13.6
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"01000001011001001100110011001100"), -- 9.2 + 5.1 = 14.3
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"10111101110011001100110011000000"), -- -5 + 4.9 = -0.0999999
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000000100101100110011001100110"), -- 4 + -8.7 = -4.7
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000001010100011001100110011001"), -- -4.7 + -8.4 = -13.1
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000000000000000000000000000010"), -- -7.1 + 9.1 = 2
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"00111111010011001100110011001100"), -- -0.1 + 0.9 = 0.8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000001001100110011001100110011"), -- 3.6 + 7.6 = 11.2
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000001100110011001100110011"), -- 0.8 + -3.6 = -2.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000001000101100110011001100110"), -- -2.8 + -6.6 = -9.4
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000000000011001100110011001101"), -- -3.5 + 1.3 = -2.2
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000001001001001100110011001101"), -- -7.8 + -2.5 = -10.3
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000001000111100110011001100110"), -- -4.9 + -5 = -9.9
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000001001100011001100110011010"), -- 5.5 + 5.6 = 11.1
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000011000000000000000000000"), -- -5.8 + 9.3 = 3.5
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111000110011001100110011010"), -- -2.2 + 1.6 = -0.6
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000000101001100110011001100111"), -- -0.6 + 5.8 = 5.2
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"10111110110011001100110011001100"), -- -2.3 + 1.9 = -0.4
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000000111000000000000000000000"), -- 2.4 + 4.6 = 7
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000001000100011001100110011010"), -- 0.5 + -9.6 = -9.1
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"00111110100110011001100110010000"), -- 4.7 + -4.4 = 0.3
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"11000000010001100110011001100111"), -- -5.3 + 2.2 = -3.1
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000000100100000000000000000000"), -- 3.8 + -8.3 = -4.5
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000010001100110011001100110"), -- -4.1 + 7.2 = 3.1
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000000001100110011001100110011"), -- 3.6 + -0.8 = 2.8
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000000100000000000000000000000"), -- 0.5 + -4.5 = -4
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"00111111001100110011001100110011"), -- 0.7 + -0 = 0.7
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000000011001100110011001101"), -- -0 + -2.2 = -2.2
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000001110011001100110011010"), -- 1.1 + 1.8 = 2.9
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"10111111101001100110011001101000"), -- 6 + -7.3 = -1.3
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000000111001100110011001100110"), -- 0.3 + -7.5 = -7.2
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"10111111011001100110011001100100"), -- 1.2 + -2.1 = -0.9
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"00111111101100110011001100110100"), -- 8.5 + -7.1 = 1.4
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000001010000000000000000000000"), -- 9 + 3 = 12
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"01000000110111001100110011001100"), -- 1.8 + 5.1 = 6.9
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101100000000000000000000"), -- -3.9 + -1.6 = -5.5
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"10111111110110011001100110011000"), -- 5.4 + -7.1 = -1.7
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000110001100110011001100110"), -- -3.4 + -2.8 = -6.2
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001010110110011001100110011"), -- -5.5 + -8.2 = -13.7
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000000110000110011001100110011"), -- 2.4 + -8.5 = -6.1
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001010110000000000000000000"), -- -4.6 + -8.9 = -13.5
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000001001111100110011001100110"), -- 7.8 + 4.1 = 11.9
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001010000011001100110011010"), -- 7.9 + 4.2 = 12.1
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000000101100110011001100110011"), -- -2.3 + -3.3 = -5.6
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"11000000001000000000000000000001"), -- -6.3 + 3.8 = -2.5
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"00111101110011001100110011000000"), -- 5.4 + -5.3 = 0.0999999
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"10111111100000000000000000000000"), -- 4.9 + -5.9 = -1
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001000011001100110011001100"), -- -3.1 + -5.7 = -8.8
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111111100110011001100110100"), -- 4.3 + -2.4 = 1.9
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"01000001010100011001100110011010"), -- 6.2 + 6.9 = 13.1
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001000110000000000000000000"), -- -1 + -8.5 = -9.5
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000000100010011001100110011010"), -- -1.3 + 5.6 = 4.3
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000000101010011001100110011001"), -- 3.4 + -8.7 = -5.3
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000001100101011001100110011010"), -- 9.5 + 9.2 = 18.7
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000001001010000000000000000000"), -- -4.9 + -5.6 = -10.5
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"10111111101001100110011001101000"), -- 4.6 + -5.9 = -1.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000000110011001100110011001100"), -- -3.5 + 9.9 = 6.4
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000001001100110011001100110011"), -- 2.5 + 8.7 = 11.2
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"01000001001010000000000000000000"), -- 2.2 + 8.3 = 10.5
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000000000110011001100110011010"), -- -2.7 + 0.3 = -2.4
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001001111100110011001100110"), -- -4.4 + -7.5 = -11.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"01000001000010011001100110011010"), -- -0 + 8.6 = 8.6
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000001100000001100110011001101"), -- 7.9 + 8.2 = 16.1
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111011001100110011001101", b"11000000111011001100110011001101"), -- 0 + -7.4 = -7.4
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"10111111011001100110011001110000"), -- 8.7 + -9.6 = -0.900001
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"10111111000000000000000000000000"), -- -8.9 + 8.4 = -0.5
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000001000100000000000000000000"), -- 9.3 + -0.3 = 9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000001010010110011001100110100"), -- 2.9 + 9.8 = 12.7
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000101100000000000000000000"), -- -5.3 + -0.2 = -5.5
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000001010000011001100110011010"), -- 6.7 + 5.4 = 12.1
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000000111000000000000000000000"), -- -2.7 + 9.7 = 7
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"00111111010011001100110011010000"), -- -7.8 + 8.6 = 0.8
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"11000001001001001100110011001101"), -- -6 + -4.3 = -10.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000111000110011001100110011"), -- -3.6 + -3.5 = -7.1
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"00111111111001100110011001101000"), -- 7.4 + -5.6 = 1.8
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000000111100110011001100110100"), -- 4.3 + 3.3 = 7.6
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000000111111001100110011001101"), -- 0.1 + 7.8 = 7.9
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001011110000000000000000000"), -- -7 + -8.5 = -15.5
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"01000000011001100110011001100110"), -- 7.5 + -3.9 = 3.6
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"01000001000011001100110011001101"), -- 1.3 + 7.5 = 8.8
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000100000000000000000000", b"00111111111001100110011001101000"), -- -7.2 + 9 = 1.8
	(b"11000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"11000000010000000000000000000000"), -- -8.8 + 5.8 = -3
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000101011001100110011001101"), -- 2.7 + 2.7 = 5.4
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000001001000011001100110011010"), -- -4.3 + -5.8 = -10.1
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000100111001100110011001100"), -- -1.3 + -3.6 = -4.9
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000001000100110011001100110011"), -- 9.5 + -0.3 = 9.2
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001001010011001100110011010"), -- 3.4 + 7.2 = 10.6
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000001000010000000000000000000"), -- -6.4 + -2.1 = -8.5
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000111100000000000000000000"), -- 5 + 2.5 = 7.5
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000001010010110011001100110100"), -- -4.1 + -8.6 = -12.7
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000001001000000000000000000000"), -- -0.7 + -9.3 = -10
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000000101000000000000000000000"), -- 3.3 + 1.7 = 5
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000001010000011001100110011010"), -- 5.6 + 6.5 = 12.1
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000000011110011001100110011010"), -- -0.5 + -3.4 = -3.9
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000100000000000000000000", b"00111111010011001100110011010000"), -- -8.2 + 9 = 0.8
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000001010111001100110011001100"), -- -8.2 + -5.6 = -13.8
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"10111101110011001100110011000000"), -- -3 + 2.9 = -0.0999999
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"11000000111100110011001100110010"), -- -9.4 + 1.8 = -7.6
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000001001110000000000000000000"), -- -9.6 + -1.9 = -11.5
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"10111110010011001100110011010000"), -- 1.8 + -2 = -0.2
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000001000011001100110011001101"), -- 5.3 + 3.5 = 8.8
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"01000000001001100110011001100110"), -- 6.5 + -3.9 = 2.6
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"00111111110110011001100110011100"), -- -3.1 + 4.8 = 1.7
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000101110011001100110011010"), -- -4.6 + -1.2 = -5.8
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000001000100000000000000000000"), -- -5.5 + -3.5 = -9
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"01000000001000000000000000000000"), -- -3.4 + 5.9 = 2.5
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"00111110110011001100110011010000"), -- -7.5 + 7.9 = 0.4
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001000000110011001100110011"), -- -4.5 + -3.7 = -8.2
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"11000000100100000000000000000000"), -- -6.3 + 1.8 = -4.5
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000000100000110011001100110100"), -- 3.8 + -7.9 = -4.1
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001100010000000000000000000"), -- -8.3 + -8.7 = -17
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000001001010110011001100110100"), -- 3.9 + 6.8 = 10.7
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000100010011001100110011010"), -- -1.1 + -3.2 = -4.3
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000001001111001100110011001101"), -- 6.5 + 5.3 = 11.8
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000000100010011001100110011010"), -- -3.1 + 7.4 = 4.3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000100010011001100110011001"), -- 0.7 + 3.6 = 4.3
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000001010100000000000000000000"), -- 3.2 + 9.8 = 13
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001100101100110011001100110"), -- 9.1 + 9.7 = 18.8
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"01000001001011001100110011001101"), -- 5.8 + 5 = 10.8
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000000000100110011001100110010"), -- 4.3 + -6.6 = -2.3
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000001001010000000000000000000"), -- 4.9 + 5.6 = 10.5
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"01000000011000000000000000000000"), -- -3.1 + 6.6 = 3.5
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000101110011001100110011010"), -- 7.3 + -1.5 = 5.8
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000001000001100110011001100110"), -- -1 + 9.4 = 8.4
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"00111110010011001100110011000000"), -- -9.1 + 9.3 = 0.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000000111000110011001100110100"), -- -0.2 + 7.3 = 7.1
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"00111110100110011001100110011000"), -- 3.5 + -3.2 = 0.3
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"01000000100111001100110011001101"), -- 7.9 + -3 = 4.9
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001010111100110011001100110"), -- 4.4 + 9.5 = 13.9
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"10111110111111111111111111110000"), -- 7.9 + -8.4 = -0.5
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"01000001010110011001100110011010"), -- 6.7 + 6.9 = 13.6
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000001001110000000000000000000"), -- -8 + -3.5 = -11.5
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000000010001100110011001100110"), -- -2.6 + 5.7 = 3.1
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"11000000101011001100110011001110"), -- 3.7 + -9.1 = -5.4
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000000011100110011001100110100"), -- -2.5 + 6.3 = 3.8
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"01000000011011001100110011001100"), -- 7.1 + -3.4 = 3.7
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000000100010011001100110011010"), -- -3.3 + 7.6 = 4.3
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"01000000110100000000000000000000"), -- 1.4 + 5.1 = 6.5
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000001010011001100110011001101"), -- 6.5 + 6.3 = 12.8
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"10111111001100110011001100111000"), -- 7.1 + -7.8 = -0.7
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000110100110011001100110100"), -- -1.8 + -4.8 = -6.6
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000000100101100110011001100110"), -- -0.5 + 5.2 = 4.7
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000001000110000000000000000000"), -- -4.5 + -5 = -9.5
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"10111111110000000000000000000000"), -- 3 + -4.5 = -1.5
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"11000000000000000000000000000000"), -- -8.7 + 6.7 = -2
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001000110110011001100110011"), -- -1.5 + -8.2 = -9.7
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000000111000000000000000000000"), -- -0.7 + -6.3 = -7
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000000111000110011001100110100"), -- 1.7 + -8.8 = -7.1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"01000000101000110011001100110011"), -- 0.6 + 4.5 = 5.1
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"10111111001100110011001100110000"), -- 8 + -8.7 = -0.7
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000000101000000000000000000000"), -- -3.5 + 8.5 = 5
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001011100110011001100110011"), -- -7 + -8.2 = -15.2
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000001001000011001100110011001"), -- -8.9 + -1.2 = -10.1
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"11000000111110011001100110011010"), -- -3.2 + -4.6 = -7.8
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000000011001100110011001100110"), -- -2.5 + 6.1 = 3.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"00111110110011001100110011001100"), -- 1.5 + -1.1 = 0.4
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"00111101110011001100110011000000"), -- 7.9 + -7.8 = 0.0999999
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000001010010011001100110011001"), -- 9.9 + 2.7 = 12.6
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001001010011001100110011010"), -- -5.3 + -5.3 = -10.6
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000001000000011001100110011010"), -- -3.9 + -4.2 = -8.1
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000001011100110011001100110100"), -- -6.6 + -8.6 = -15.2
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"01000000000110011001100110011010"), -- -4.5 + 6.9 = 2.4
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000000101101100110011001100111"), -- 3.1 + -8.8 = -5.7
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"11000000010100110011001100110100"), -- -9 + 5.7 = -3.3
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000000100111111111111111111111"), -- -4.4 + 9.4 = 5
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001011010011001100110011010"), -- 5 + 9.6 = 14.6
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000000000011001100110011001100"), -- 7.7 + -9.9 = -2.2
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000010001100110011001100110"), -- -1.9 + -1.2 = -3.1
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001011100011001100110011010"), -- -5.6 + -9.5 = -15.1
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001100101000000000000000000"), -- 9 + 9.5 = 18.5
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"11000000110111111111111111111111"), -- -9.9 + 2.9 = -7
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000110111001100110011001101"), -- 5.9 + 1 = 6.9
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000010110011001100110011010"), -- 1.8 + 1.6 = 3.4
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"), -- -7.7 + 7.7 = 0
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"01000000101100000000000000000000"), -- 8 + -2.5 = 5.5
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"01000001010110110011001100110100"), -- 7.3 + 6.4 = 13.7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000000110011001100110011001"), -- -2.8 + 0.4 = -2.4
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"11000000001011001100110011001100"), -- -6.6 + 3.9 = -2.7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"10111111111100110011001100110010"), -- 3.7 + -5.6 = -1.9
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000000100110011001100110100"), -- -4.9 + 2.6 = -2.3
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111111100110011001100110011001"), -- -1.1 + 2.3 = 1.2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000001000001001100110011001101"), -- -2.5 + -5.8 = -8.3
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000111011001100110011001101"), -- 3.7 + 3.7 = 7.4
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"10111111011001100110011001101000"), -- -6.1 + 5.2 = -0.9
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001001111100110011001100110"), -- -3.2 + -8.7 = -11.9
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"11000001011111001100110011001100"), -- -8.9 + -6.9 = -15.8
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"00111111111001100110011001101000"), -- -5.7 + 7.5 = 1.8
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000000111000110011001100110010"), -- -1.3 + 8.4 = 7.1
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000001000010011001100110011010"), -- 1.5 + 7.1 = 8.6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000000101000110011001100110011"), -- 0.8 + -5.9 = -5.1
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000110101100110011001100110"), -- -6 + -0.7 = -6.7
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000000101000110011001100110011"), -- 2.4 + -7.5 = -5.1
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"01000001011000011001100110011010"), -- 9.1 + 5 = 14.1
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001010000011001100110011010"), -- -6.4 + -5.7 = -12.1
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001011001100110011001100110"), -- 4.9 + 9.5 = 14.4
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000010100110011001100110011"), -- -3.1 + -0.2 = -3.3
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000001000001001100110011001100"), -- -5.7 + -2.6 = -8.3
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001010000110011001100110100"), -- -4.3 + -7.9 = -12.2
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001001110110011001100110011"), -- 2 + 9.7 = 11.7
	(b"11000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000001011000110011001100110011"), -- -8.4 + -5.8 = -14.2
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"11000001010000011001100110011010"), -- -7.5 + -4.6 = -12.1
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111101110011001100110011100000"), -- -2.9 + 2.8 = -0.1
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001010110000000000000000000"), -- 3.8 + 9.7 = 13.5
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000000111000110011001100110011"), -- 0.6 + 6.5 = 7.1
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000000110011001100110011001"), -- 0.1 + 2.3 = 2.4
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000001001110000000000000000000"), -- 3.1 + 8.4 = 11.5
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"10111111110110011001100110011100"), -- -5.3 + 3.6 = -1.7
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"10111111110011001100110011001100"), -- 4.1 + -5.7 = -1.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"01000001000001001100110011001101"), -- 3.5 + 4.8 = 8.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"10111111100011001100110011001110"), -- 2.8 + -3.9 = -1.1
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"10111110110011001100110011001000"), -- 3.7 + -4.1 = -0.4
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000001100000110011001100110100"), -- 9.6 + 6.8 = 16.4
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000000110100110011001100110011"), -- -1.9 + 8.5 = 6.6
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"10111111001100110011001100110010"), -- 1.1 + -1.8 = -0.7
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"11000000111100110011001100110011"), -- -9.7 + 2.1 = -7.6
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000001001011001100110011001101"), -- -9.5 + -1.3 = -10.8
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000100001100110011001100111"), -- -5.1 + 9.3 = 4.2
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"01000000101010011001100110011001"), -- 7.2 + -1.9 = 5.3
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000000111011001100110011001101"), -- -6.5 + -0.9 = -7.4
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"00111111111001100110011001100000"), -- -8.1 + 9.9 = 1.8
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000001000110011001100110011010"), -- 8.8 + 0.8 = 9.6
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000101110011001100110011010"), -- 6.8 + -1 = 5.8
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001011001100110011001100110"), -- 8.3 + 6.1 = 14.4
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"10111111111100110011001100110100"), -- -9.5 + 7.6 = -1.9
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001001001001100110011001101"), -- -6.6 + -3.7 = -10.3
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000001001110110011001100110100"), -- 6.8 + 4.9 = 11.7
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"01000000101010011001100110011001"), -- 8.4 + -3.1 = 5.3
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000100000000000000000000", b"01000001100101000000000000000000"), -- 9.5 + 9 = 18.5
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000100010011001100110011010"), -- 4.9 + -0.6 = 4.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"11000001000000011001100110011010"), -- -1 + -7.1 = -8.1
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001100100001100110011001100"), -- -8.7 + -9.4 = -18.1
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000100000110011001100110100"), -- -5.3 + 1.2 = -4.1
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"00111111100110011001100110011100"), -- 8.8 + -7.6 = 1.2
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"00111111110000000000000000000000"), -- 9.8 + -8.3 = 1.5
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"01000000011000000000000000000000"), -- 5.4 + -1.9 = 3.5
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000000000000000000000000000000"), -- 7.8 + -9.8 = -2
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"01000001000100011001100110011010"), -- 4.6 + 4.5 = 9.1
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000001000001100110011001100110"), -- -2.5 + -5.9 = -8.4
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"01000000010011001100110011001101"), -- 5.5 + -2.3 = 3.2
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"00111111011001100110011001100100"), -- 4.2 + -3.3 = 0.9
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000001011110110011001100110011"), -- -9.2 + -6.5 = -15.7
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111111110000000000000000000000"), -- -2.1 + 3.6 = 1.5
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"01000000100000110011001100110100"), -- -1.8 + 5.9 = 4.1
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"01000000100100000000000000000000"), -- 6.5 + -2 = 4.5
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"01000000110110011001100110011001"), -- 8.4 + -1.6 = 6.8
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000001100001001100110011001101"), -- 7.9 + 8.7 = 16.6
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100010011001100110011010", b"01000001000000011001100110011010"), -- 3.8 + 4.3 = 8.1
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"01000000111100110011001100110011"), -- 9 + -1.4 = 7.6
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"00111111001100110011001100110000"), -- -8.2 + 8.9 = 0.7
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"10111111001100110011001100110000"), -- -5.6 + 4.9 = -0.7
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000001001000011001100110011001"), -- 8.9 + 1.2 = 10.1
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000000100111111111111111111111"), -- -3.4 + 8.4 = 5
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000001100001011001100110011010"), -- 9.4 + 7.3 = 16.7
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000100100110011001100110011"), -- 2.3 + 2.3 = 4.6
	(b"01000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100011001100110011001101", b"01000001000110011001100110011010"), -- 5.2 + 4.4 = 9.6
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000000011011001100110011001100"), -- 6.2 + -9.9 = -3.7
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001010000110011001100110011"), -- -7.7 + -4.5 = -12.2
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001100010110011001100110011"), -- -9.9 + -7.5 = -17.4
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"10111110110011001100110011010000"), -- -8.3 + 7.9 = -0.4
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111011001100110011001101", b"10111111111001100110011001101000"), -- 5.6 + -7.4 = -1.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"10111111101111111111111111111110"), -- 3.7 + -5.2 = -1.5
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"11000001000110011001100110011010"), -- -2.5 + -7.1 = -9.6
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001010100000000000000000000"), -- 6 + 7 = 13
	(b"11000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"), -- -4.8 + 4.8 = 0
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"10111111110110011001100110011010"), -- -2.9 + 1.2 = -1.7
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000010011001100110011001100"), -- -1 + 4.2 = 3.2
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"10111111101001100110011001100111"), -- 1.9 + -3.2 = -1.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000001010000011001100110011010"), -- 2.8 + 9.3 = 12.1
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000001000000000000000000000000"), -- -4.1 + -3.9 = -8
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000001000010000000000000000000"), -- -4.3 + -4.2 = -8.5
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000001000000000000000000000000"), -- 7.6 + 0.4 = 8
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000001000000011001100110011010"), -- 4.3 + 3.8 = 8.1
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"), -- 7.4 + -7.4 = 0
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000001011110000000000000000000"), -- -8.9 + -6.6 = -15.5
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001001101100110011001100110"), -- -6.1 + -5.3 = -11.4
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000101111001100110011001101"), -- 6 + -0.1 = 5.9
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000000010011001100110011001100"), -- -2.4 + 5.6 = 3.2
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"00111111110110011001100110011000"), -- 8.4 + -6.7 = 1.7
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000001000100000000000000000000"), -- -0.3 + 9.3 = 9
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000001000100000000000000000000"), -- 0.6 + -9.6 = -9
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000101010011001100110011010"), -- 4.5 + 0.8 = 5.3
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000000110000000000000000000000"), -- -1.1 + -4.9 = -6
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001100010001100110011001101"), -- 7.6 + 9.5 = 17.1
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"10111111001100110011001100111000"), -- -7.4 + 6.7 = -0.7
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000100100110011001100110100"), -- 0.2 + -4.8 = -4.6
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000001010000000000000000000000"), -- -8.1 + -3.9 = -12
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001010110011001100110011001"), -- -4.2 + -9.4 = -13.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111100000000000000000000000"), -- 2 + -1 = 1
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000111101100110011001100110"), -- -6.7 + -1 = -7.7
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001000111100110011001100110"), -- -5 + -4.9 = -9.9
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000100011001100110011001101"), -- -2.2 + -2.2 = -4.4
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"01000000001011001100110011001110"), -- -4.2 + 6.9 = 2.7
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000001000101001100110011001101"), -- -3.5 + -5.8 = -9.3
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000001010010110011001100110100"), -- 7.8 + 4.9 = 12.7
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000100010011001100110011010"), -- -2.1 + -2.2 = -4.3
	(b"01000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"01000000100100110011001100110011"), -- 8.2 + -3.6 = 4.6
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000001000110110011001100110011"), -- -2.5 + -7.2 = -9.7
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000001011001100110011001101"), -- 2.3 + 0.4 = 2.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000100101100110011001100110"), -- 2.6 + 2.1 = 4.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000000111111001100110011001101"), -- 2.6 + 5.3 = 7.9
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000000011100110011001100110010"), -- -5.9 + 9.7 = 3.8
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"00111111000110011001100110010000"), -- 8.9 + -8.3 = 0.599999
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"11000000000100110011001100110100"), -- -3.4 + 1.1 = -2.3
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000001010111001100110011001101"), -- -7 + -6.8 = -13.8
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000001001010110011001100110011"), -- 7.1 + 3.6 = 10.7
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000000111011001100110011001110"), -- -1.7 + 9.1 = 7.4
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000111101100110011001100110"), -- 5 + 2.7 = 7.7
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"01000000110011001100110011001101"), -- 8.8 + -2.4 = 6.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001000000011001100110011010"), -- -0 + -8.1 = -8.1
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000000101001100110011001100110"), -- -6.5 + 1.3 = -5.2
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000000111101100110011001100110"), -- 8.5 + -0.8 = 7.7
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000101000000000000000000000"), -- -2.1 + -2.9 = -5
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"10111101110011001100110011001100"), -- 0.3 + -0.4 = -0.1
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001100010100110011001100110"), -- -8.6 + -8.7 = -17.3
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"01000001000010110011001100110011"), -- 4 + 4.7 = 8.7
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"00111110100110011001100110010000"), -- 4.7 + -4.4 = 0.3
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000001100100000000000000000000"), -- -9.2 + -8.8 = -18
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"00111111110110011001100110011010"), -- -1.3 + 3 = 1.7
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000001000100000000000000000000"), -- -9.7 + 0.7 = -9
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"10111111110011001100110011001100"), -- -7.9 + 6.3 = -1.6
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000000010001100110011001100111"), -- 2.2 + -5.3 = -3.1
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000001001100000000000000000000"), -- -8.6 + -2.4 = -11
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"00111111010011001100110011010000"), -- -4.1 + 4.9 = 0.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000001000000011001100110011010"), -- -0 + 8.1 = 8.1
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000001001000110011001100110100"), -- -8.1 + -2.1 = -10.2
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"01000000000110011001100110011010"), -- 7.9 + -5.5 = 2.4
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001010100110011001100110011"), -- -4.5 + -8.7 = -13.2
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001011010110011001100110011"), -- -6.7 + -8 = -14.7
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100010011001100110011010", b"01000001000100011001100110011010"), -- 4.8 + 4.3 = 9.1
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000000111100110011001100110011"), -- 0.9 + -8.5 = -7.6
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000000100000110011001100110011"), -- -4.7 + 0.6 = -4.1
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001010110000000000000000000"), -- 7.4 + 6.1 = 13.5
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000101000110011001100110011"), -- 2.3 + 2.8 = 5.1
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000001001010011001100110011010"), -- -8.5 + -2.1 = -10.6
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000001011111100110011001100110"), -- 7.4 + 8.5 = 15.9
	(b"01000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"00111111100011001100110011001100"), -- 5.7 + -4.6 = 1.1
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000000101110011001100110011010"), -- 1.2 + 4.6 = 5.8
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000001100010110011001100110100"), -- -8.1 + -9.3 = -17.4
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"10111111010011001100110011010000"), -- -9.1 + 8.3 = -0.8
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101100000000000000000000", b"01000001001010000000000000000000"), -- 5 + 5.5 = 10.5
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000101110011001100110011001"), -- 0.9 + -6.7 = -5.8
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101011001100110011001100"), -- -2.8 + -2.6 = -5.4
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001000100011001100110011001"), -- -0.9 + -8.2 = -9.1
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000001011001100110011001101"), -- -1 + -1.7 = -2.7
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"11000000100000000000000000000000"), -- -7.1 + 3.1 = -4
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000101110011001100110011001"), -- 1.6 + 4.2 = 5.8
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001010001100110011001100110"), -- -8.7 + -3.7 = -12.4
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001001110011001100110011010"), -- 2 + 9.6 = 11.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001001010000000000000000000"), -- 3.3 + 7.2 = 10.5
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100011001100110011001101", b"11000000010110011001100110011010"), -- -7.8 + 4.4 = -3.4
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000001000010011001100110011010"), -- -0 + -8.6 = -8.6
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000001000000011001100110011010"), -- -6.8 + -1.3 = -8.1
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001010011100110011001100110"), -- 3.2 + 9.7 = 12.9
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000000110000000000000000000000"), -- 0.3 + 5.7 = 6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001001001001100110011001100"), -- -1.4 + -8.9 = -10.3
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000000111100110011001100110011"), -- 0.9 + -8.5 = -7.6
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"11000000101110011001100110011010"), -- 1.2 + -7 = -5.8
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000000101111001100110011001101"), -- -0.9 + -5 = -5.9
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"10111111000000000000000000000000"), -- 0 + -0.5 = -0.5
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"00111111101001100110011001101000"), -- -7.5 + 8.8 = 1.3
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"11000000100010011001100110011010"), -- -9.5 + 5.2 = -4.3
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000001001111001100110011001101"), -- -8.5 + -3.3 = -11.8
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000000110100110011001100110100"), -- -1.3 + -5.3 = -6.6
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000000100100110011001100110011"), -- -0.1 + -4.5 = -4.6
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001010100000000000000000000"), -- -4.1 + -8.9 = -13
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000000101000000000000000000000"), -- 0.2 + -5.2 = -5
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000000011001100110011001100111"), -- -0.4 + -3.2 = -3.6
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000000111111001100110011001101"), -- 0.4 + -8.3 = -7.9
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000101100110011001100110011"), -- 6 + -0.4 = 5.6
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000001010110000000000000000000"), -- 5.6 + 7.9 = 13.5
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000000111011001100110011001101"), -- -0.8 + -6.6 = -7.4
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111101110011001100110011001101"), -- -0.1 + 0.2 = 0.1
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111111100110011001100110011"), -- 1.9 + -3.8 = -1.9
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001001011001100110011001100"), -- -1.4 + -9.4 = -10.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001100110011001100110011"), -- -0 + -2.8 = -2.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000000011110011001100110011010"), -- 3.9 + -0 = 3.9
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000001001000110011001100110011"), -- 8 + 2.2 = 10.2
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001001000000000000000000000"), -- -3.7 + -6.3 = -10
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000100011001100110011001101"), -- 0.5 + 3.9 = 4.4
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000001011000000000000000000000"), -- 7.8 + 6.2 = 14
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000110000000000000000000000"), -- 3 + 3 = 6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"10111111011001100110011001100100"), -- 2.7 + -3.6 = -0.9
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"00111111101001100110011001101000"), -- -8 + 9.3 = 1.3
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001000100110011001100110011"), -- -4.7 + -4.5 = -9.2
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000001011001100110011001101"), -- 4.4 + -1.7 = 2.7
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"01000000010100110011001100110010"), -- 8.7 + -5.4 = 3.3
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000000100100000000000000000001"), -- 4.1 + -8.6 = -4.5
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000000100111001100110011001100"), -- 4.5 + -9.4 = -4.9
	(b"01000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"01000000001100110011001100110100"), -- 8.6 + -5.8 = 2.8
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000000011110011001100110011010"), -- -4.9 + 8.8 = 3.9
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000000010000000000000000000000"), -- 4.5 + -7.5 = -3
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"10111111111001100110011001101000"), -- 2.5 + -4.3 = -1.8
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001000011001100110011001101"), -- -5.1 + -3.7 = -8.8
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000001001001001100110011001101"), -- 9.6 + 0.7 = 10.3
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000001010011100110011001100110"), -- 9.3 + 3.6 = 12.9
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"11000000100001100110011001100110"), -- -6.5 + 2.3 = -4.2
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000001001000000000000000000000"), -- -1.7 + -8.3 = -10
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101100000000000000000000", b"01000001010100110011001100110011"), -- 7.7 + 5.5 = 13.2
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000001011000110011001100110100"), -- -4.4 + -9.8 = -14.2
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000000100110011001100110011"), -- 0.4 + 1.9 = 2.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"), -- 0.6 + -0.6 = 0
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000001000110110011001100110011"), -- -7.4 + -2.3 = -9.7
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"01000000101101100110011001100110"), -- 0.6 + 5.1 = 5.7
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001010010000000000000000000"), -- -7.3 + -5.2 = -12.5
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"01000000100111001100110011001100"), -- 7.6 + -2.7 = 4.9
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"10111111000000000000000000000000"), -- 0.5 + -1 = -0.5
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"11000001100010011001100110011010"), -- -8.1 + -9.1 = -17.2
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"00111111100000000000000000000000"), -- -8.6 + 9.6 = 1
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"), -- -4.7 + 4.7 = 0
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"10111110110011001100110011010000"), -- -6.1 + 5.7 = -0.4
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111100110011001100110011010"), -- -0.4 + -0.8 = -1.2
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"10111111011001100110011001100000"), -- 5.3 + -6.2 = -0.9
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000001001010110011001100110011"), -- -7.7 + -3 = -10.7
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000111111001100110011001101"), -- -7.1 + -0.8 = -7.9
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001000100000000000000000000"), -- 4.8 + 4.2 = 9
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000101010011001100110011010"), -- -1.6 + -3.7 = -5.3
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000001011001100110011001100"), -- 0.4 + -3.1 = -2.7
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000000010011001100110011001110"), -- -4.7 + 7.9 = 3.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"00111111100000000000000000000000"), -- 3.2 + -2.2 = 1
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000010001100110011001100110"), -- -0.6 + 3.7 = 3.1
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000001010000011001100110011010"), -- 5.4 + 6.7 = 12.1
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001011101001100110011001101"), -- 8.1 + 7.2 = 15.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"00111111110011001100110011001101"), -- -0.6 + 2.2 = 1.6
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"01000000010110011001100110011010"), -- 6.5 + -3.1 = 3.4
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"11000001000000011001100110011001"), -- -8.9 + 0.8 = -8.1
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"10111101110011001100110100000000"), -- -5.8 + 5.7 = -0.1
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001011110000000000000000000"), -- 8.5 + 7 = 15.5
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001011100000000000000000000"), -- 5.3 + 9.7 = 15
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000001000011001100110011001101"), -- -7.9 + -0.9 = -8.8
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"01000000100001100110011001100110"), -- 6 + -1.8 = 4.2
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000001000000110011001100110011"), -- -0 + 8.2 = 8.2
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"00111101110011001100110011000000"), -- -2.2 + 2.3 = 0.0999999
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111001100110011001100110011"), -- 0.5 + 0.2 = 0.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"11000001001101100110011001100110"), -- -3.6 + -7.8 = -11.4
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"11000001010100110011001100110100"), -- -5.4 + -7.8 = -13.2
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000100010011001100110011010"), -- 1.2 + 3.1 = 4.3
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001000000000000000000000000"), -- -2.8 + -5.2 = -8
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001010000011001100110011010"), -- -4.6 + -7.5 = -12.1
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11000000000100110011001100110011"), -- -2.3 + 0 = -2.3
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000001001010011001100110011001"), -- -9.2 + -1.4 = -10.6
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000000100000000000000000000000"), -- -3.9 + 7.9 = 4
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000001100000011001100110011010"), -- -7 + -9.2 = -16.2
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"00111111110110011001100110011100"), -- 6.3 + -4.6 = 1.7
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"10111110100110011001100110100000"), -- -7.3 + 7 = -0.3
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"11000000100011001100110011001100"), -- -7.2 + 2.8 = -4.4
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000001000000011001100110011001"), -- -1.9 + -6.2 = -8.1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000000100110011001100110011010"), -- 0.6 + -5.4 = -4.8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000000011001100110011001101"), -- -0.3 + 2.5 = 2.2
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"10111110010011001100110011100000"), -- -5.8 + 5.6 = -0.2
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001011100011001100110011001"), -- -9.4 + -5.7 = -15.1
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001100001110011001100110011"), -- -7.5 + -9.4 = -16.9
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"10111111110110011001100110011100"), -- 4.2 + -5.9 = -1.7
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"10111111111100110011001100110100"), -- 4.7 + -6.6 = -1.9
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000000111111001100110011001101"), -- -1.9 + -6 = -7.9
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000001000101001100110011001100"), -- -8.9 + -0.4 = -9.3
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000001100000100110011001100110"), -- -8.6 + -7.7 = -16.3
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001010000011001100110011010"), -- -7.2 + -4.9 = -12.1
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000001000101001100110011001101"), -- 0.2 + 9.1 = 9.3
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000001011011100110011001100110"), -- -8.9 + -6 = -14.9
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000111100110011001100110100"), -- 4.8 + 2.8 = 7.6
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000001100010011001100110011010"), -- 9.8 + 7.4 = 17.2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000000101001100110011001100110"), -- -2.5 + 7.7 = 5.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000111000000000000000000000"), -- -0.2 + -6.8 = -7
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"01000000011000000000000000000001"), -- 7.3 + -3.8 = 3.5
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"10111111111001100110011001100110"), -- 1.7 + -3.5 = -1.8
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"00111111111001100110011001100100"), -- -4.9 + 6.7 = 1.8
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"01000000100000000000000000000000"), -- 9.3 + -5.3 = 4
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000001010110110011001100110100"), -- -8.1 + -5.6 = -13.7
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000000111000000000000000000000"), -- -1.3 + -5.7 = -7
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000001100001100110011001100110"), -- -8.2 + -8.6 = -16.8
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001100001000000000000000000"), -- -9 + -7.5 = -16.5
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000001010000110011001100110100"), -- 4.4 + 7.8 = 12.2
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000101101100110011001100110"), -- 6.7 + -1 = 5.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000000110110011001100110011010"), -- 2.2 + 4.6 = 6.8
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000000111110011001100110011001"), -- 2.6 + 5.2 = 7.8
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"11000000110001100110011001100110"), -- -1.1 + -5.1 = -6.2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000000111101100110011001100110"), -- -1.2 + 8.9 = 7.7
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000001100101000000000000000000"), -- 9.3 + 9.2 = 18.5
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000001001100110011001100110100"), -- -9.1 + -2.1 = -11.2
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000010001100110011001101000"), -- -6.2 + 9.3 = 3.1
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000000101110011001100110011010"), -- -0 + 5.8 = 5.8
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000001000000110011001100110011"), -- 0 + 8.2 = 8.2
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"00111111000110011001100110100000"), -- 9.1 + -8.5 = 0.6
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"11000000011100110011001100110100"), -- -6.3 + 2.5 = -3.8
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000010011001100110011001101"), -- 3 + 0.2 = 3.2
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"00111111001100110011001100111000"), -- 7.9 + -7.2 = 0.7
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"01000000111010011001100110011001"), -- 0.7 + 6.6 = 7.3
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001010100011001100110011001"), -- 8.9 + 4.2 = 13.1
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"11000000100011001100110011001101"), -- -7.8 + 3.4 = -4.4
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"11000000001011001100110011001101"), -- -6 + 3.3 = -2.7
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000101010011001100110011001"), -- 4.7 + 0.6 = 5.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"11000000100100000000000000000000"), -- 0.6 + -5.1 = -4.5
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000100111001100110011001101"), -- 3.9 + 1 = 4.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000100010011001100110011010"), -- -3.5 + -0.8 = -4.3
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"01000001100011110011001100110100"), -- 9.3 + 8.6 = 17.9
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"01000000100100000000000000000000"), -- 6.4 + -1.9 = 4.5
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"01000000100001100110011001100110"), -- 9.7 + -5.5 = 4.2
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001010101100110011001100110"), -- -4.4 + -9 = -13.4
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001011000011001100110011001"), -- 9.9 + 4.2 = 14.1
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001100010001100110011001101"), -- 7.4 + 9.7 = 17.1
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000011000000000000000000000"), -- 1.7 + 1.8 = 3.5
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111101001100110011001100110"), -- 1.5 + -2.8 = -1.3
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"00111111100110011001100110011000"), -- 7.5 + -6.3 = 1.2
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001100101011001100110011010"), -- 9 + 9.7 = 18.7
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000001000100000000000000000000"), -- 9.2 + -0.2 = 9
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001001000011001100110011001"), -- 0.4 + 9.7 = 10.1
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"11000001000001100110011001100111"), -- -0.6 + -7.8 = -8.4
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"01000000100000110011001100110100"), -- 9.8 + -5.7 = 4.1
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000111100110011001100110011"), -- -6.9 + -0.7 = -7.6
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000001000010000000000000000000"), -- -7.6 + -0.9 = -8.5
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000000001000000000000000000000"), -- 1.6 + -4.1 = -2.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000000110110011001100110011010"), -- 1.9 + 4.9 = 6.8
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"10111111001100110011001100110000"), -- -6.1 + 5.4 = -0.7
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000001100001000000000000000000"), -- 8.3 + 8.2 = 16.5
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000100000000000000000000000"), -- -1.8 + -2.2 = -4
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000000101101100110011001100110"), -- -3 + 8.7 = 5.7
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001000010011001100110011010"), -- -0.1 + -8.5 = -8.6
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000000111101100110011001100110"), -- 2 + 5.7 = 7.7
	(b"11000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"11000000001100110011001100110100"), -- -9.8 + 7 = -2.8
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000001000100110011001100110011"), -- 5.1 + 4.1 = 9.2
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"11000000111100110011001100110011"), -- -8.7 + 1.1 = -7.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000000101001100110011001100110"), -- 3.5 + -8.7 = -5.2
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000001000000000000000000000000"), -- 1.3 + -9.3 = -8
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001011000011001100110011010"), -- -9.6 + -4.5 = -14.1
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"00111111110011001100110011010000"), -- -6.7 + 8.3 = 1.6
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"01000001001000110011001100110011"), -- 5.5 + 4.7 = 10.2
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000001001000011001100110011010"), -- 3.4 + 6.7 = 10.1
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"11000000010100110011001100110011"), -- -3 + -0.3 = -3.3
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000001000110000000000000000000"), -- 1.7 + 7.8 = 9.5
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000001000010110011001100110011"), -- 6.2 + 2.5 = 8.7
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001100100110011001100110011"), -- -9.5 + -8.9 = -18.4
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111100011001100110011001101"), -- -0.5 + 1.6 = 1.1
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000001001110110011001100110100"), -- 8.8 + 2.9 = 11.7
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000001000110011001100110011010"), -- -5.4 + -4.2 = -9.6
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000000100000110011001100110100"), -- -1.2 + 5.3 = 4.1
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000001010010011001100110011010"), -- 4.1 + 8.5 = 12.6
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"11000001010011100110011001100110"), -- -7.8 + -5.1 = -12.9
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000000100001100110011001100110"), -- -2 + 6.2 = 4.2
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101100000000000000000000", b"01000000110000000000000000000000"), -- 0.5 + 5.5 = 6
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"01000001010110110011001100110011"), -- 7.7 + 6 = 13.7
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"11000000101101100110011001100110"), -- -1.7 + -4 = -5.7
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000000101111001100110011001101"), -- -1.5 + -4.4 = -5.9
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"00111110110011001100110011100000"), -- -8.9 + 9.3 = 0.400001
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000001000101001100110011001101"), -- -5.4 + -3.9 = -9.3
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000000111111001100110011001101"), -- 8.8 + -0.9 = 7.9
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000001100001001100110011001101"), -- -7.4 + -9.2 = -16.6
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000001100000000000000000000000"), -- -8.7 + -7.3 = -16
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000001000000110011001100110011"), -- -1.1 + 9.3 = 8.2
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"10111110010011001100110011000000"), -- 6.9 + -7.1 = -0.2
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000000111010011001100110011001"), -- 2.1 + 5.2 = 7.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000111010011001100110011001"), -- -0.6 + -6.7 = -7.3
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001000100011001100110011010"), -- -0.5 + 9.6 = 9.1
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000111000110011001100110100"), -- -3.4 + -3.7 = -7.1
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"01000000011100110011001100110100"), -- -3.1 + 6.9 = 3.8
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"01000000100000000000000000000000"), -- 7.4 + -3.4 = 4
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"11000000011011001100110011001110"), -- -9.6 + 5.9 = -3.7
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000001010110011001100110011010"), -- -7.1 + -6.5 = -13.6
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"11000000010110011001100110011010"), -- -5.8 + 2.4 = -3.4
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"10111111111100110011001100110011"), -- -3 + 1.1 = -1.9
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001000010011001100110011001"), -- 0.1 + -8.7 = -8.6
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000100000000000000000000", b"01000001000100000000000000000000"), -- -0 + 9 = 9
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000001001100110011001100110100"), -- -2.4 + -8.8 = -11.2
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000001000110011001100110011010"), -- -9.1 + -0.5 = -9.6
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000000000110011001100110011010"), -- 4.9 + -7.3 = -2.4
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000001110011001100110011001"), -- 0.7 + -3.6 = -2.9
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000001001100000000000000000000"), -- 8.3 + 2.7 = 11
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000001000101100110011001100110"), -- -7.2 + -2.2 = -9.4
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000001000001001100110011001101"), -- 9.1 + -0.8 = 8.3
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000001001010110011001100110100"), -- -8.6 + -2.1 = -10.7
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"00111111010011001100110011001000"), -- 4.7 + -3.9 = 0.8
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"00111111101001100110011001101000"), -- -5.5 + 6.8 = 1.3
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"11000000000110011001100110011010"), -- -4 + 1.6 = -2.4
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"11000000000000000000000000000010"), -- -9.6 + 7.6 = -2
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000001100110011001100110100"), -- 4 + -6.8 = -2.8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000000010000000000000000000000"), -- 3.6 + -6.6 = -3
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001001110011001100110011001"), -- -2.2 + -9.4 = -11.6
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000010111111111111111111111"), -- -3.7 + 7.2 = 3.5
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000001100001110011001100110011"), -- 9.8 + 7.1 = 16.9
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000010100110011001100110100"), -- 3.9 + -0.6 = 3.3
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000100101100110011001100110"), -- -4.2 + -0.5 = -4.7
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000101001100110011001100110"), -- 4.2 + 1 = 5.2
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111101001100110011001100110"), -- 1.4 + -0.1 = 1.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000000001110011001100110011010"), -- -1.2 + -1.7 = -2.9
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000001100100011001100110011010"), -- 8.3 + 9.9 = 18.2
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"11000000110000110011001100110011"), -- -9.5 + 3.4 = -6.1
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001100000011001100110011010"), -- 9 + 7.2 = 16.2
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000100100000000000000000000"), -- 4.1 + 0.4 = 4.5
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000001010110110011001100110011"), -- -9.9 + -3.8 = -13.7
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"11000000101010011001100110011001"), -- -7.2 + 1.9 = -5.3
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000010011001100110011001100"), -- -1.8 + -1.4 = -3.2
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"11000000001100110011001100110100"), -- -8.1 + 5.3 = -2.8
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001000000110011001100110011"), -- -0.2 + -8 = -8.2
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000000000001100110011001100111"), -- 1.8 + -3.9 = -2.1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000000000001100110011001100110"), -- 2.1 + -4.2 = -2.1
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000111111001100110011001100"), -- 6.7 + 1.2 = 7.9
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000000101010011001100110011010"), -- -1.5 + 6.8 = 5.3
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000001011101100110011001100110"), -- -8.9 + -6.5 = -15.4
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"11000000101100110011001100110011"), -- -6.6 + 1 = -5.6
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000000111100000000000000000000"), -- -2.2 + 9.7 = 7.5
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000010000000000000000000000"), -- 1.1 + 1.9 = 3
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"01000000010001100110011001100110"), -- 7.6 + -4.5 = 3.1
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001011100110011001100110011"), -- -7.2 + -8 = -15.2
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"00111110100110011001100110100000"), -- 9.3 + -9 = 0.3
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"00111111110110011001100110011001"), -- -1.6 + 3.3 = 1.7
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000111100110011001100110011"), -- -6.6 + -1 = -7.6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000000111100110011001100110011"), -- -1.4 + -6.2 = -7.6
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"11000000100000000000000000000000"), -- 3.1 + -7.1 = -4
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"01000000100011001100110011001101"), -- 3.3 + 1.1 = 4.4
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"00111111000000000000000000000000"), -- 6.8 + -6.3 = 0.5
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000110000110011001100110011"), -- 3.6 + 2.5 = 6.1
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000001010101100110011001100110"), -- 4.9 + 8.5 = 13.4
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000001000100000000000000000000"), -- 8.9 + 0.1 = 9
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000111010011001100110011010"), -- 9 + -1.7 = 7.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"00111101110011001100110011010000"), -- -1 + 1.1 = 0.1
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000101100000000000000000000"), -- 5.1 + 0.4 = 5.5
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000000001100110011001100111"), -- 1.7 + 0.4 = 2.1
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"11000000111100000000000000000000"), -- -9.5 + 2 = -7.5
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001001011100110011001100110"), -- -2.7 + -8.2 = -10.9
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000000000110011001100110011001"), -- -3.7 + 6.1 = 2.4
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000001001110011001100110011010"), -- -6.6 + -5 = -11.6
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"00111110010011001100110011100000"), -- 4.8 + -4.6 = 0.2
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"11000000101100000000000000000000"), -- -1.5 + -4 = -5.5
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000000110010011001100110011010"), -- 5.1 + 1.2 = 6.3
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000001010101100110011001100110"), -- -6.6 + -6.8 = -13.4
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"00111110100110011001100110010000"), -- -5.3 + 5.6 = 0.3
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"00111111100011001100110011001100"), -- 7.9 + -6.8 = 1.1
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"11000000010001100110011001100111"), -- -5.9 + 2.8 = -3.1
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001011010110011001100110011"), -- -6.7 + -8 = -14.7
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000110111001100110011001100"), -- -0.3 + 7.2 = 6.9
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"01000000011001100110011001100111"), -- 7.4 + -3.8 = 3.6
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000110000000000000000000000"), -- -4.5 + -1.5 = -6
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"10111110010011001100110011010000"), -- -3.9 + 3.7 = -0.2
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000001000111001100110011001101"), -- 1.1 + 8.7 = 9.8
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000011000000000000000000000"), -- 0.5 + 3 = 3.5
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"11000001011101100110011001100110"), -- -8.3 + -7.1 = -15.4
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"01000000111100000000000000000000"), -- 8.8 + -1.3 = 7.5
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000001100110011001100110011"), -- 2.1 + 0.7 = 2.8
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"01000001010001100110011001100110"), -- 5.8 + 6.6 = 12.4
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000001001001100110011001100110"), -- 4.2 + 6.2 = 10.4
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000000111000110011001100110010"), -- -2.3 + 9.4 = 7.1
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"10111111011001100110011001101000"), -- -8.3 + 7.4 = -0.9
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"10111111010011001100110011001100"), -- 2 + -2.8 = -0.8
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"11000000001011001100110011001100"), -- -9 + 6.3 = -2.7
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000100011001100110011001100"), -- -5.6 + 1.2 = -4.4
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"00111111110110011001100110011000"), -- 6.2 + -4.5 = 1.7
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000001000100110011001100110011"), -- -1.9 + -7.3 = -9.2
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000000101100110011001100110100"), -- -0.2 + 5.8 = 5.6
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000010100110011001100110100"), -- 4.3 + -1 = 3.3
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001001001100110011001100110"), -- -4.7 + -5.7 = -10.4
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000010011001100110011001101"), -- -3.7 + 0.5 = -3.2
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"10111111100110011001100110011000"), -- 5 + -6.2 = -1.2
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000001010011001100110011001100"), -- 8.7 + 4.1 = 12.8
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000001010000011001100110011010"), -- 6.7 + 5.4 = 12.1
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"10111110100110011001100110100000"), -- 7.8 + -8.1 = -0.3
	(b"01000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"00111111001100110011001100110000"), -- 8.2 + -7.5 = 0.7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000000001000000000000000000000"), -- -3.6 + 6.1 = 2.5
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001011110000000000000000000"), -- -7.4 + -8.1 = -15.5
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"01000000101110011001100110011010"), -- 7.9 + -2.1 = 5.8
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000101110011001100110011010"), -- -3.3 + -2.5 = -5.8
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001010000110011001100110100"), -- -7.3 + -4.9 = -12.2
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000001011000110011001100110011"), -- 9 + 5.2 = 14.2
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"00111111110011001100110011001100"), -- 9.2 + -7.6 = 1.6
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"00111111011001100110011001101000"), -- 7.9 + -7 = 0.9
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000000111001100110011001100110"), -- 0.1 + 7.1 = 7.2
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100101100110011001100110", b"01000000010001100110011001101000"), -- 7.8 + -4.7 = 3.1
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000000111100000000000000000000"), -- -3.3 + -4.2 = -7.5
	(b"01000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000001001100110011001100110011"), -- 6.6 + 4.6 = 11.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000000101010011001100110011010"), -- -0.9 + -4.4 = -5.3
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000000110000110011001100110011"), -- -0.4 + 6.5 = 6.1
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000111100000000000000000000"), -- -5.2 + -2.3 = -7.5
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"), -- 0.7 + -0.7 = 0
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000111101100110011001100111"), -- -8.1 + 0.4 = -7.7
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001011111001100110011001101"), -- -7.7 + -8.1 = -15.8
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000000011110011001100110011010"), -- 1 + 2.9 = 3.9
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000001000110011001100110011010"), -- -6.3 + -3.3 = -9.6
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000001001101001100110011001100"), -- -7.7 + -3.6 = -11.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000000111100000000000000000000"), -- -1.2 + -6.3 = -7.5
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000001100001100110011001100110"), -- -6.9 + -9.9 = -16.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000000110101100110011001100110"), -- -0 + 6.7 = 6.7
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111111111100110011001100110011"), -- -1.9 + 3.8 = 1.9
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000001000000000000000000000000"), -- 7.8 + 0.2 = 8
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"01000000101110011001100110011001"), -- 0.7 + 5.1 = 5.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"10111111110110011001100110011000"), -- 3.9 + -5.6 = -1.7
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"01000000100001100110011001100111"), -- 7.8 + -3.6 = 4.2
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"01000000100100110011001100110011"), -- 9.7 + -5.1 = 4.6
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000001001000110011001100110011"), -- 9.5 + 0.7 = 10.2
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001011101100110011001100110"), -- -5.7 + -9.7 = -15.4
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"11000001001110000000000000000000"), -- -5.4 + -6.1 = -11.5
	(b"01000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"01000000100000110011001100110011"), -- 5.7 + -1.6 = 4.1
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001000100011001100110011001"), -- 0.3 + -9.4 = -9.1
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"10111111110000000000000000000000"), -- -0.7 + -0.8 = -1.5
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"01000000000100110011001100110100"), -- -6 + 8.3 = 2.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000000101101100110011001100111"), -- -0.6 + 6.3 = 5.7
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"01000000101000000000000000000000"), -- 0.3 + 4.7 = 5
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"10111111110110011001100110011000"), -- -5.6 + 3.9 = -1.7
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000100110011001100110011010"), -- 5.5 + -0.7 = 4.8
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"01000000010011001100110011001110"), -- 8.1 + -4.9 = 3.2
	(b"01000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"01000000101000000000000000000001"), -- 8.6 + -3.6 = 5
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000111000110011001100110100"), -- -8.3 + 1.2 = -7.1
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000001010110011001100110011010"), -- 6 + 7.6 = 13.6
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000000001001100110011001100110"), -- 0.2 + -2.8 = -2.6
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000011110011001100110011010"), -- -0.9 + -3 = -3.9
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000001000010011001100110011010"), -- 7.9 + 0.7 = 8.6
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000100000110011001100110100"), -- 2.7 + -6.8 = -4.1
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"11000000011000000000000000000000"), -- -6 + 2.5 = -3.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000000100110011001100110011"), -- 1.9 + 0.4 = 2.3
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"01000000100100110011001100110011"), -- -1.4 + 6 = 4.6
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"00111111101001100110011001100110"), -- -1.3 + 2.6 = 1.3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000001010010000000000000000000"), -- 2.6 + 9.9 = 12.5
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001001011001100110011001101"), -- -1.8 + -9 = -10.8
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000111001100110011001100111"), -- -5.3 + -1.9 = -7.2
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"11000001000000000000000000000000"), -- -9.6 + 1.6 = -8
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"11000000101100110011001100110010"), -- -9.4 + 3.8 = -5.6
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000001000001100110011001100110"), -- 1.5 + -9.9 = -8.4
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"11000000110010011001100110011010"), -- -1.7 + -4.6 = -6.3
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001010101001100110011001100"), -- -5.7 + -7.6 = -13.3
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000000010011001100110011001100"), -- 4.1 + -0.9 = 3.2
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"01000000000110011001100110011010"), -- 7.4 + -5 = 2.4
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000000100110011001100110011001"), -- 4.6 + -9.4 = -4.8
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000000100111001100110011001101"), -- -4.1 + -0.8 = -4.9
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000001001011001100110011001101"), -- -7.6 + -3.2 = -10.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000101010011001100110011001"), -- 1.4 + -6.7 = -5.3
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111111101001100110011001100110"), -- 3.1 + -1.8 = 1.3
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001001100110011001100110011"), -- 4.2 + 7 = 11.2
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"00111111100000000000000000000000"), -- 9.5 + -8.5 = 1
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000001010101001100110011001100"), -- 9.2 + 4.1 = 13.3
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001001100011001100110011010"), -- 6.9 + 4.2 = 11.1
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000101111001100110011001101"), -- 2.5 + 3.4 = 5.9
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000000111001100110011001100110"), -- 4.1 + 3.1 = 7.2
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000000111010011001100110011001"), -- 2.6 + -9.9 = -7.3
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"00111111111100110011001100110011"), -- -0 + 1.9 = 1.9
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000001010011001100110011001101"), -- 3.2 + 9.6 = 12.8
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000100100110011001100110011"), -- 2 + 2.6 = 4.6
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"01000001001100011001100110011010"), -- 6.1 + 5 = 11.1
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"00111111000000000000000000000000"), -- 6.8 + -6.3 = 0.5
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000001001100110011001100111"), -- 2.2 + -4.8 = -2.6
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"), -- -2.4 + 2.4 = 0
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000000100001100110011001100111"), -- 0.2 + -4.4 = -4.2
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000000101100000000000000000000"), -- 0.1 + 5.4 = 5.5
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001011100110011001100110011"), -- -6.7 + -8.5 = -15.2
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111111000110011001100110011001"), -- -1.4 + 0.8 = -0.6
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000001001001001100110011001100"), -- -9.4 + -0.9 = -10.3
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000000100101100110011001100111"), -- 0.6 + -5.3 = -4.7
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000000110011001100110011001100"), -- -2 + 8.4 = 6.4
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"00111111011001100110011001100000"), -- 7.2 + -6.3 = 0.9
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"01000000001000000000000000000000"), -- 7.3 + -4.8 = 2.5
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"10111111100110011001100110011001"), -- -2.8 + 1.6 = -1.2
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000001001011001100110011001100"), -- 5.6 + 5.2 = 10.8
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"11000000101011001100110011001110"), -- -9.6 + 4.2 = -5.4
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"11000001000000000000000000000000"), -- -9.6 + 1.6 = -8
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001001111001100110011001100"), -- 7.6 + 4.2 = 11.8
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000110100110011001100110011"), -- 7 + -0.4 = 6.6
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"00111101110011001100110011000000"), -- 3.6 + -3.5 = 0.0999999
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000001011110110011001100110011"), -- 6.8 + 8.9 = 15.7
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000000111000110011001100110011"), -- -1.4 + -5.7 = -7.1
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000001001010110011001100110011"), -- 3.1 + 7.6 = 10.7
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"10111111000110011001100110011000"), -- 5.8 + -6.4 = -0.6
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000100001100110011001100111"), -- 4.8 + -0.6 = 4.2
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000001001011100110011001100110"), -- 7.4 + 3.5 = 10.9
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"11000001011100110011001100110011"), -- -9.7 + -5.5 = -15.2
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000000111011001100110011001101"), -- 8 + -0.6 = 7.4
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"11000000101010011001100110011010"), -- -8.6 + 3.3 = -5.3
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000001010000110011001100110100"), -- -9.1 + -3.1 = -12.2
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"01000000101000000000000000000000"), -- -1.6 + 6.6 = 5
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"10111110100110011001100110100000"), -- 8.9 + -9.2 = -0.3
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"10111111101100110011001100110100"), -- 3.6 + -5 = -1.4
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"00111111100110011001100110011010"), -- 1 + 0.2 = 1.2
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"11000000110111001100110011001100"), -- -4.2 + -2.7 = -6.9
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000001010000011001100110011010"), -- 9.1 + 3 = 12.1
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000001000111001100110011001100"), -- 9.9 + -0.1 = 9.8
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000001100001100110011001100110"), -- 7 + 9.8 = 16.8
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001011110110011001100110011"), -- -6.7 + -9 = -15.7
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"11000001011100000000000000000000"), -- -8.1 + -6.9 = -15
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"00111111110110011001100110011001"), -- 1.8 + -0.1 = 1.7
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000001100111011001100110011010"), -- 9.8 + 9.9 = 19.7
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001010110110011001100110011"), -- -8.5 + -5.2 = -13.7
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000011001100110011001100110"), -- -1.4 + -2.2 = -3.6
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"11000000010100110011001100110100"), -- -7.5 + 4.2 = -3.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001001100110011001100110"), -- 2.8 + -0.2 = 2.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"10111111101001100110011001101000"), -- 3.5 + -4.8 = -1.3
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000011001100110011001100110"), -- -6.2 + 2.6 = -3.6
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000010000000000000000000000"), -- 3.3 + -0.3 = 3
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000000000011001100110011001110"), -- -3.1 + 5.3 = 2.2
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000101111001100110011001101"), -- -3.4 + 9.3 = 5.9
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000001000010110011001100110011"), -- -1 + -7.7 = -8.7
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100011001100110011001101", b"11000000101100110011001100110011"), -- -6.7 + 1.1 = -5.6
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000100000110011001100110011"), -- -3.1 + 7.2 = 4.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111111001100110011001100111"), -- -1.2 + -0.6 = -1.8
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000010001100110011001100110"), -- -1 + -2.1 = -3.1
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000001010100110011001100110100"), -- -7.4 + -5.8 = -13.2
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000000100110011001100110011001"), -- -2.9 + 7.7 = 4.8
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000101100000000000000000000"), -- -3.8 + 9.3 = 5.5
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000110001100110011001100110"), -- 3.2 + 3 = 6.2
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000001000011100110011001100110"), -- 9 + -0.1 = 8.9
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000000100000110011001100110100"), -- 5.5 + -9.6 = -4.1
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"00111110010011001100110100000000"), -- 9.1 + -8.9 = 0.200001
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000001000010000000000000000000"), -- -4.9 + -3.6 = -8.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000000101100000000000000000000"), -- 0.4 + -5.9 = -5.5
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"01000001011110000000000000000000"), -- 9.6 + 5.9 = 15.5
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000011000000000000000000000"), -- 1.4 + 2.1 = 3.5
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"00111111100011001100110011001100"), -- 7.1 + -6 = 1.1
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000001010111100110011001100110"), -- -7.1 + -6.8 = -13.9
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000001001010011001100110011010"), -- -5.6 + -5 = -10.6
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000000100010011001100110011010"), -- -3.8 + -0.5 = -4.3
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000001001101100110011001100110"), -- -1.5 + -9.9 = -11.4
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"10111101110011001100110100000000"), -- -8.3 + 8.2 = -0.1
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000111000110011001100110011"), -- -7.1 + -0 = -7.1
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001011010110011001100110011"), -- -6.2 + -8.5 = -14.7
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000000110000000000000000000000"), -- 3.7 + -9.7 = -6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000000000001100110011001100110"), -- 0.8 + 1.3 = 2.1
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"11000000010011001100110011001100"), -- -9.9 + 6.7 = -3.2
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001100010000000000000000000"), -- -7.5 + -9.5 = -17
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000000111011001100110011001100"), -- -2.2 + -5.2 = -7.4
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000000000110011001100110011010"), -- -7.4 + 9.8 = 2.4
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"00111111001100110011001100110000"), -- -5.5 + 6.2 = 0.7
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"10111111011001100110011001100000"), -- 6.8 + -7.7 = -0.9
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000000110000000000000000000000"), -- -3.7 + 9.7 = 6
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"00111111000110011001100110011000"), -- 7 + -6.4 = 0.6
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"10111111111100110011001100110100"), -- 4.7 + -6.6 = -1.9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000000110010011001100110011001"), -- 2.9 + -9.2 = -6.3
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000000001110011001100110011010"), -- 6.1 + -9 = -2.9
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000001000001100110011001100110"), -- -9.7 + 1.3 = -8.4
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"01000000011001100110011001100100"), -- 8.4 + -4.8 = 3.6
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"01000001001100000000000000000000"), -- 6.3 + 4.7 = 11
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000000011100110011001100110010"), -- 6.1 + -9.9 = -3.8
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000000111000110011001100110011"), -- 1.4 + -8.5 = -7.1
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000000100101100110011001100110"), -- -4.7 + 9.4 = 4.7
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000001000010110011001100110100"), -- 9.6 + -0.9 = 8.7
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000000101000000000000000000001"), -- 4.6 + -9.6 = -5
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000001011001001100110011001100"), -- -5.4 + -8.9 = -14.3
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"01000001000100110011001100110011"), -- 9.8 + -0.6 = 9.2
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000000110000000000000000000000"), -- 1.9 + 4.1 = 6
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"00111101110011001100110011000000"), -- 6 + -5.9 = 0.0999999
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"10111111100000000000000000000000"), -- -8.7 + 7.7 = -1
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"11000000101111001100110011001101"), -- -0.4 + -5.5 = -5.9
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000001010100110011001100110011"), -- -6.5 + -6.7 = -13.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111100011001100110011001101"), -- -0.5 + 1.6 = 1.1
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001000101100110011001100110"), -- 3.3 + 6.1 = 9.4
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000001001011100110011001100110"), -- 9.5 + 1.4 = 10.9
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000100000000000000000000000"), -- 2.4 + 1.6 = 4
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000001000110000000000000000000"), -- 9.8 + -0.3 = 9.5
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000000100111001100110011001101"), -- -0.8 + -4.1 = -4.9
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001001111100110011001100110"), -- 5.8 + 6.1 = 11.9
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000011110011001100110011010"), -- 2.5 + 1.4 = 3.9
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"10111110100110011001100110000000"), -- 8.1 + -8.4 = -0.299999
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000000110011001100110011010"), -- -5 + 2.6 = -2.4
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000110000110011001100110011"), -- -1.1 + 7.2 = 6.1
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"01000001000011001100110011001101"), -- 8.5 + 0.3 = 8.8
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001011011100110011001100111"), -- -6.8 + -8.1 = -14.9
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000000101100000000000000000000"), -- 1 + -6.5 = -5.5
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001011101100110011001100110"), -- -5.9 + -9.5 = -15.4
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"01000000001011001100110011001100"), -- 7.1 + -4.4 = 2.7
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"11000001001010011001100110011010"), -- -5.5 + -5.1 = -10.6
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"01000000100000000000000000000000"), -- 7.8 + -3.8 = 4
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000001001100000000000000000000"), -- 2.9 + 8.1 = 11
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001010010000000000000000000"), -- -8 + -4.5 = -12.5
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001000010000000000000000000"), -- -0.3 + -8.2 = -8.5
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001000110000000000000000000"), -- -1.9 + -7.6 = -9.5
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000000110010011001100110011010"), -- 3.5 + -9.8 = -6.3
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000110000000000000000000000"), -- 3.7 + 2.3 = 6
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001000011100110011001100110"), -- 1.7 + 7.2 = 8.9
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000000110000000000000000000000"), -- 1.3 + -7.3 = -6
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000001000010110011001100110011"), -- -3.1 + -5.6 = -8.7
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000000101111001100110011001100"), -- 3.8 + -9.7 = -5.9
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000110100110011001100110100"), -- -2.7 + 9.3 = 6.6
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000101000110011001100110011"), -- 5.4 + -0.3 = 5.1
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000001000000000000000000000"), -- 3.6 + -1.1 = 2.5
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000001000011001100110011001101"), -- 8.3 + 0.5 = 8.8
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"11000000001011001100110011001100"), -- -8.9 + 6.2 = -2.7
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"11000000100000000000000000000000"), -- -8.2 + 4.2 = -4
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000000000100110011001100110100"), -- 2.1 + -4.4 = -2.3
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"11000000011001100110011001100110"), -- -7.5 + 3.9 = -3.6
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"11000000001000000000000000000000"), -- -9.5 + 7 = -2.5
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"11000000100111001100110011001100"), -- -8.7 + 3.8 = -4.9
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"10111111111100110011001100110000"), -- 8 + -9.9 = -1.9
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000001000000011001100110011001"), -- 8.4 + -0.3 = 8.1
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000001011000000000000000000000"), -- 6.7 + 7.3 = 14
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001000001001100110011001101"), -- -0.7 + -7.6 = -8.3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000001000100011001100110011010"), -- 2.6 + 6.5 = 9.1
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000100101100110011001100110"), -- -2.9 + -1.8 = -4.7
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000000101100000000000000000000"), -- 7.2 + -1.7 = 5.5
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000000001000000000000000000000"), -- -2.1 + -0.4 = -2.5
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"11000000100011001100110011001110"), -- -9.1 + 4.7 = -4.4
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001011111100110011001100111"), -- -9.6 + -6.3 = -15.9
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"10111101110011001100110011000000"), -- -3.8 + 3.7 = -0.0999999
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"01000000000001100110011001100110"), -- 5 + -2.9 = 2.1
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000001010100011001100110011010"), -- 6 + 7.1 = 13.1
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110110011001100110011010"), -- -3.9 + -2.9 = -6.8
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000100100000000000000000000"), -- 2.2 + -6.7 = -4.5
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000001001101100110011001100110"), -- -7.9 + -3.5 = -11.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000000101101100110011001100110"), -- 0 + -5.7 = -5.7
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000001011010000000000000000000"), -- -6.1 + -8.4 = -14.5
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001110011001100110011010", b"01000001000101100110011001100110"), -- 6.5 + 2.9 = 9.4
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"10111111100110011001100110011001"), -- -1.3 + 0.1 = -1.2
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"01000001011100011001100110011010"), -- 8.7 + 6.4 = 15.1
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000001100001110011001100110011"), -- -8.5 + -8.4 = -16.9
	(b"01000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"01000000100011001100110011001110"), -- 8.6 + -4.2 = 4.4
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"00111111110110011001100110011000"), -- 7.2 + -5.5 = 1.7
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000001010000000000000000000000"), -- -4.3 + -7.7 = -12
	(b"11000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001011001001100110011001101"), -- -9.8 + -4.5 = -14.3
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000001001001001100110011001101"), -- 7.8 + 2.5 = 10.3
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000001000011001100110011001101"), -- 9.7 + -0.9 = 8.8
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"01000000010001100110011001100111"), -- 5.3 + -2.2 = 3.1
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"10111111111001100110011001101000"), -- 7.7 + -9.5 = -1.8
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"11000001000000110011001100110011"), -- -9.7 + 1.5 = -8.2
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000001001100110011001100110011"), -- 7.5 + 3.7 = 11.2
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"), -- -8 + 8 = 0
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000110001100110011001100110"), -- -3.3 + -2.9 = -6.2
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"00111110110011001100110011010000"), -- 3.4 + -3 = 0.4
	(b"01000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"01000000111100110011001100110010"), -- 9.9 + -2.3 = 7.6
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000001010001001100110011001101"), -- 9.5 + 2.8 = 12.3
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"11000001000010011001100110011010"), -- -6.9 + -1.7 = -8.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000110110011001100110011010"), -- -2 + -4.8 = -6.8
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000000010110011001100110011010"), -- 3 + -6.4 = -3.4
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000001001011100110011001100110"), -- 7.6 + 3.3 = 10.9
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001001000110011001100110011"), -- -0.5 + -9.7 = -10.2
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"01000000000001100110011001100110"), -- 7.9 + -5.8 = 2.1
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000001001000011001100110011010"), -- 2.7 + 7.4 = 10.1
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"10111111000000000000000000000000"), -- 6.3 + -6.8 = -0.5
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"01000000000000000000000000000000"), -- 4.6 + -2.6 = 2
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001011100011001100110011010"), -- -5.4 + -9.7 = -15.1
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001011100000000000000000000"), -- -7.1 + -7.9 = -15
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"11000000010000000000000000000000"), -- -6.5 + 3.5 = -3
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"01000000100101100110011001100110"), -- 8.4 + -3.7 = 4.7
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001001001001100110011001100"), -- 6.1 + 4.2 = 10.3
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000000101100000000000000000000"), -- 1 + -6.5 = -5.5
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"01000000110100000000000000000000"), -- -1.5 + 8 = 6.5
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000001000110110011001100110100"), -- 0.6 + 9.1 = 9.7
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111111101001100110011001100110"), -- -4.1 + 2.8 = -1.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001000010110011001100110100"), -- -0.6 + -8.1 = -8.7
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000001000100110011001100110011"), -- 0 + 9.2 = 9.2
	(b"11000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"11000000110001100110011001100111"), -- -9.8 + 3.6 = -6.2
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"11000000101111001100110011001100"), -- -9.4 + 3.5 = -5.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000101000110011001100110011"), -- -3.5 + -1.6 = -5.1
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000001001000011001100110011010"), -- -5.7 + -4.4 = -10.1
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000000011100110011001100110100"), -- 1.1 + -4.9 = -3.8
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"11000001000100110011001100110011"), -- -3.7 + -5.5 = -9.2
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000001001110011001100110011010"), -- -9.3 + -2.3 = -11.6
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000000100111001100110011001100"), -- 1.3 + -6.2 = -4.9
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000000010011001100110011001101"), -- 1.7 + -4.9 = -3.2
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"11000001010011001100110011001101"), -- -8.6 + -4.2 = -12.8
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000001100101100110011001100110"), -- 9.1 + 9.7 = 18.8
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000000011001100110011001101"), -- 0.8 + 1.4 = 2.2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"00111111100011001100110011001101"), -- 0.7 + 0.4 = 1.1
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"01000000010000000000000000000000"), -- 7.9 + -4.9 = 3
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000110011001100110011001100"), -- 2.6 + 3.8 = 6.4
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"11000001000010000000000000000000"), -- -7.7 + -0.8 = -8.5
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"10111111111001100110011001100111"), -- -1.2 + -0.6 = -1.8
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"01000000001100110011001100110010"), -- 9.2 + -6.4 = 2.8
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000001000111001100110011001101"), -- -3.4 + -6.4 = -9.8
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001001011001100110011001101"), -- -1.1 + -9.7 = -10.8
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000001000110000000000000000000"), -- -6.4 + -3.1 = -9.5
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000000011011001100110011001100"), -- 1.1 + 2.6 = 3.7
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"00111111110000000000000000000000"), -- -7.2 + 8.7 = 1.5
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"10111101110011001100110011100000"), -- -3.4 + 3.3 = -0.1
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"10111111000110011001100110011000"), -- 3.5 + -4.1 = -0.6
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"11000000100100110011001100110100"), -- -7.8 + 3.2 = -4.6
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"11000000001110011001100110011010"), -- -6.9 + 4 = -2.9
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"11000000100010011001100110011010"), -- -9.3 + 5 = -4.3
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"01000000001011001100110011001100"), -- -5.3 + 8 = 2.7
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"01000000100100000000000000000000"), -- 6.3 + -1.8 = 4.5
	(b"11000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001001000011001100110011010"), -- -4.8 + -5.3 = -10.1
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"10111111000000000000000000000000"), -- -7.3 + 6.8 = -0.5
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000001001111100110011001100110"), -- -8.5 + -3.4 = -11.9
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"01000001100100001100110011001101"), -- 9.5 + 8.6 = 18.1
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000001011110110011001100110011"), -- 6.8 + 8.9 = 15.7
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"00111111010011001100110011001100"), -- -2.7 + 3.5 = 0.8
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"01000000001100110011001100110100"), -- 7.8 + -5 = 2.8
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"01000000000011001100110011001100"), -- 8.4 + -6.2 = 2.2
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"10111111100110011001100110011010"), -- -1 + -0.2 = -1.2
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"00111110110011001100110011010000"), -- 3 + -2.6 = 0.4
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000101011001100110011001101"), -- 2.7 + 2.7 = 5.4
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"01000000001100110011001100110011"), -- 5 + -2.2 = 2.8
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100011001100110011001101", b"01000001001010000000000000000000"), -- 6.1 + 4.4 = 10.5
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000110011001100110011001101"), -- 5.8 + 0.6 = 6.4
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000000001100110011001100110100"), -- 3.6 + -6.4 = -2.8
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"11000000010011001100110011001101"), -- -6 + 2.8 = -3.2
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000111100110011001100110011"), -- 8 + -0.4 = 7.6
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"00111110010011001100110011001100"), -- -0.3 + 0.5 = 0.2
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000100111001100110011001101"), -- 3.5 + 1.4 = 4.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000000001011001100110011001100"), -- -0.9 + -1.8 = -2.7
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000000111100000000000000000000"), -- 1.8 + -9.3 = -7.5
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000001010101001100110011001100"), -- -3.4 + -9.9 = -13.3
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000001001001001100110011001100"), -- 3.1 + 7.2 = 10.3
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"01000000100111001100110011001101"), -- 7.5 + -2.6 = 4.9
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000101001100110011001100111"), -- -7.8 + 2.6 = -5.2
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000001000011100110011001100111"), -- 7.3 + 1.6 = 8.9
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000111010011001100110011001"), -- -4.7 + -2.6 = -7.3
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"11000000110000110011001100110011"), -- -1.1 + -5 = -6.1
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000000100110011001100110011001"), -- 0.2 + 4.6 = 4.8
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000001001001001100110011001100"), -- 2.6 + 7.7 = 10.3
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"11000000010100110011001100110100"), -- -8.1 + 4.8 = -3.3
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000111010011001100110011001"), -- -6.7 + -0.6 = -7.3
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000000011110011001100110011010"), -- 4.9 + -8.8 = -3.9
	(b"01000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"01000001010100110011001100110011"), -- 5.7 + 7.5 = 13.2
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000000111011001100110011001110"), -- 0.7 + -8.1 = -7.4
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000001000100110011001100110011"), -- -3.8 + -5.4 = -9.2
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000000000000000000000000000"), -- -1 + 3 = 2
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"11000000000000000000000000000000"), -- -2.4 + 0.4 = -2
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000000100010011001100110011010"), -- 5.5 + -9.8 = -4.3
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"11000000001110011001100110011100"), -- 6.2 + -9.1 = -2.9
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"01000001011000011001100110011010"), -- 5.4 + 8.7 = 14.1
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101001100110011001100110", b"01000000101101100110011001100110"), -- 0.5 + 5.2 = 5.7
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001000111100110011001100110"), -- -5 + -4.9 = -9.9
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000000101110011001100110011010"), -- 2.5 + -8.3 = -5.8
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"11000000011001100110011001100110"), -- -5.6 + 2 = -3.6
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000001000001100110011001100110"), -- 4.6 + 3.8 = 8.4
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"01000001011110011001100110011010"), -- 7.6 + 8 = 15.6
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000111100110011001100110011"), -- -7 + -0.6 = -7.6
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001000111100110011001100110"), -- -2.3 + -7.6 = -9.9
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000100000110011001100110011"), -- 4.2 + -0.1 = 4.1
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"11000000111100110011001100110011"), -- -5.6 + -2 = -7.6
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"10111111100011001100110011001100"), -- 7.1 + -8.2 = -1.1
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"00111111111100110011001100110100"), -- 5 + -3.1 = 1.9
	(b"01000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"00111110010011001100110011000000"), -- 5.2 + -5 = 0.2
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000010001100110011001100110"), -- -0.5 + -2.6 = -3.1
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001000110110011001100110011"), -- 3.6 + 6.1 = 9.7
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000000001110011001100110011010"), -- -4.5 + 7.4 = 2.9
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000001000111001100110011001101"), -- 6 + 3.8 = 9.8
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"11000001000001001100110011001101"), -- -4 + -4.3 = -8.3
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"11000000101101100110011001100111"), -- 2.9 + -8.6 = -5.7
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"11000000101010011001100110011001"), -- -9.9 + 4.6 = -5.3
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000001001100110011001100110"), -- -1.2 + 3.8 = 2.6
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000000100011001100110011001101"), -- -3.4 + 7.8 = 4.4
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001000010000000000000000000"), -- 1.2 + -9.7 = -8.5
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000010100110011001100110100"), -- 2.9 + 0.4 = 3.3
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000001000110110011001100110011"), -- 7.6 + 2.1 = 9.7
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000001000000110011001100110011"), -- 1.4 + 6.8 = 8.2
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"00111111111001100110011001101000"), -- -3.5 + 5.3 = 1.8
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000000101111111111111111111111"), -- 2.4 + -8.4 = -6
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"10111111101100110011001100110100"), -- -8 + 6.6 = -1.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000000100100000000000000000000"), -- 3 + -7.5 = -4.5
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"11000001001001001100110011001101"), -- -6.3 + -4 = -10.3
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"10111111011001100110011001110000"), -- -8.6 + 7.7 = -0.900001
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001011101001100110011001100"), -- -6.6 + -8.7 = -15.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000000101101100110011001100110"), -- -3.5 + -2.2 = -5.7
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111110010011001100110011001100"), -- -1 + 0.8 = -0.2
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"10111111100000000000000000000001"), -- 1.9 + -2.9 = -1
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"11000000011001100110011001100110"), -- -3.5 + -0.1 = -3.6
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"10111111001100110011001100110000"), -- -4.6 + 3.9 = -0.7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"10111111100011001100110011001100"), -- -2.8 + 1.7 = -1.1
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000001001001001100110011001100"), -- -3.6 + -6.7 = -10.3
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"10111111111001100110011001100100"), -- 4.8 + -6.6 = -1.8
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000001000010011001100110011010"), -- -1.8 + -6.8 = -8.6
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000001010011001100110011001101"), -- -6 + -6.8 = -12.8
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000000011100110011001100110010"), -- -3.9 + 7.7 = 3.8
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000000110000000000000000000000"), -- 2.8 + -8.8 = -6
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000001000100011001100110011001"), -- 8.9 + 0.2 = 9.1
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000000011001100110011001101"), -- 3.2 + -1 = 2.2
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000001001110011001100110011010"), -- 5.9 + 5.7 = 11.6
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001000001001100110011001101"), -- 0.7 + -9 = -8.3
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"11000000011110011001100110011001"), -- -7.6 + 3.7 = -3.9
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000001001010000000000000000000"), -- 9 + 1.5 = 10.5
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000001010100110011001100110100"), -- 5.1 + 8.1 = 13.2
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"10111111001100110011001100111000"), -- -6.8 + 6.1 = -0.7
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"11000000111110011001100110011010"), -- -0.8 + -7 = -7.8
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"00111111011001100110011001101000"), -- -1.8 + 2.7 = 0.9
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"11000000010000000000000000000000"), -- -7.8 + 4.8 = -3
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000001100000100110011001100110"), -- -8 + -8.3 = -16.3
	(b"01000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001100000001100110011001101"), -- 6.6 + 9.5 = 16.1
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000001001000000000000000000000"), -- 2.1 + 7.9 = 10
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000000011011001100110011001101"), -- -1.2 + 4.9 = 3.7
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"01000000101000110011001100110100"), -- 5.8 + -0.7 = 5.1
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000001100000110011001100110011"), -- 8 + 8.4 = 16.4
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"11000000110001100110011001100110"), -- -7.9 + 1.7 = -6.2
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"00111111100110011001100110011100"), -- 7.9 + -6.7 = 1.2
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000001001000011001100110011010"), -- 9.3 + 0.8 = 10.1
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000010000000000000000000", b"01000001001101100110011001100110"), -- 2.9 + 8.5 = 11.4
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000110110011001100110011010"), -- 4.3 + 2.5 = 6.8
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"11000000111111001100110011001100"), -- -1.8 + -6.1 = -7.9
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000000001100110011001100110100"), -- 3.9 + -1.1 = 2.8
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"11000000100010011001100110011010"), -- -7.9 + 3.6 = -4.3
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000001000001001100110011001101"), -- 7.9 + 0.4 = 8.3
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001010101001100110011001101"), -- -8 + -5.3 = -13.3
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000000100000000000000000000000"), -- 3.6 + -7.6 = -4
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000110001100110011001100111"), -- 5.4 + 0.8 = 6.2
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"11000001000111100110011001100110"), -- -9.9 + 0 = -9.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000001100110011001100110011"), -- -3.5 + 0.7 = -2.8
	(b"01000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"01000000010000000000000000000000"), -- 9.3 + -6.3 = 3
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001011010000000000000000000"), -- -6.6 + -7.9 = -14.5
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"10111111010011001100110011001100"), -- -4.6 + 3.8 = -0.8
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000011001100110011001100110"), -- 2.7 + 0.9 = 3.6
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000001001011100110011001100110"), -- -4.4 + -6.5 = -10.9
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001010011100110011001100110"), -- -9.2 + -3.7 = -12.9
	(b"11000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"11000001000011100110011001100111"), -- -9.8 + 0.9 = -8.9
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"01000001001010011001100110011010"), -- 4.2 + 6.4 = 10.6
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000001010111100110011001100110"), -- 6.5 + 7.4 = 13.9
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000001010100011001100110011010"), -- -5.9 + -7.2 = -13.1
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001011011100110011001100111"), -- -6.8 + -8.1 = -14.9
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000010011001100110011010", b"10111111100110011001100110011100"), -- 7.4 + -8.6 = -1.2
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000000000100110011001100110010"), -- 7.6 + -9.9 = -2.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000001100110011001100110011"), -- -1 + 3.8 = 2.8
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"01000001011000000000000000000000"), -- 7.6 + 6.4 = 14
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001010000110011001100110100"), -- -6.9 + -5.3 = -12.2
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000000111001100110011001100110"), -- 0.8 + -8 = -7.2
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000000000110011001100110011010"), -- 5.5 + -7.9 = -2.4
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000001001010000000000000000000"), -- 1.3 + 9.2 = 10.5
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"00111111100000000000000000000000"), -- 2.3 + -1.3 = 1
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000001000100110011001100110100"), -- -5.3 + -3.9 = -9.2
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"00111111100000000000000000000000"), -- 7.2 + -6.2 = 1
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"10111111011001100110011001100000"), -- 8.8 + -9.7 = -0.9
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000101001100110011001100110"), -- 4.5 + 0.7 = 5.2
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"11000000100100110011001100110011"), -- -6.7 + 2.1 = -4.6
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000001000001001100110011001101"), -- -7.7 + -0.6 = -8.3
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000000111000000000000000000000"), -- -0.9 + 7.9 = 7
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001000100011001100110011010"), -- -2.8 + -6.3 = -9.1
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000000111000000000000000000000"), -- 2.3 + -9.3 = -7
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"00111111100000000000000000000000"), -- -8.7 + 9.7 = 1
	(b"11000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"10111110110011001100110011010000"), -- -3 + 2.6 = -0.4
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111101100110011001100110", b"01000001100000110011001100110011"), -- 8.7 + 7.7 = 16.4
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000001010000000000000000000000"), -- 8.8 + 3.2 = 12
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000000000000000000000000000000"), -- -0 + 2 = 2
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001100010011001100110011010"), -- -9.7 + -7.5 = -17.2
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000001011101001100110011001100"), -- 5.9 + 9.4 = 15.3
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000000100001100110011001100110"), -- 4.2 + 0 = 4.2
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000001001010011001100110011010"), -- -2.9 + -7.7 = -10.6
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000000001100110011001100110"), -- -4.7 + 2.6 = -2.1
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000000110000110011001100110011"), -- 1.1 + -7.2 = -6.1
	(b"01000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"00111111101001100110011001101000"), -- 7.9 + -6.6 = 1.3
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000010110011001100110011001"), -- -0.3 + -3.1 = -3.4
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"01000001000101001100110011001101"), -- 4.8 + 4.5 = 9.3
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"01000000001011001100110011001101"), -- 5.5 + -2.8 = 2.7
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"01000000101010011001100110011001"), -- 8.7 + -3.4 = 5.3
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000001100000001100110011001100"), -- 6.2 + 9.9 = 16.1
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000000100000000000000000000000"), -- -4.2 + 8.2 = 4
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000001011011001100110011001101"), -- 7.4 + 7.4 = 14.8
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000010000000000000000000000"), -- -5.6 + 2.6 = -3
	(b"11000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"00111111101001100110011001100100"), -- -4.8 + 6.1 = 1.3
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000001010010000000000000000000"), -- 4.4 + 8.1 = 12.5
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001000010000000000000000000"), -- -0.5 + -8 = -8.5
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"01000000100101100110011001100110"), -- 0.9 + 3.8 = 4.7
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"00111111101001100110011001100100"), -- 6.2 + -4.9 = 1.3
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000000100011001100110011001100"), -- 2.8 + -7.2 = -4.4
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000000100101100110011001100111"), -- 3.4 + -8.1 = -4.7
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000000111011001100110011001101"), -- 0.3 + 7.1 = 7.4
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000000110111001100110011001100"), -- -3.3 + -3.6 = -6.9
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000000011011001100110011001100"), -- 5.3 + -9 = -3.7
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"01000000100110011001100110011010"), -- 9.1 + -4.3 = 4.8
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"00000000000000000000000000000000", b"01000000101110011001100110011010"), -- 5.8 + 0 = 5.8
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"00111111001100110011001100110000"), -- -3.4 + 4.1 = 0.7
	(b"11000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000001100000000000000000000000"), -- -9.8 + -6.2 = -16
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101001100110011001101", b"01000000110100110011001100110100"), -- -2.7 + 9.3 = 6.6
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"01000001000111100110011001100110"), -- 7.5 + 2.4 = 9.9
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000001011000000000000000000000"), -- 7.3 + 6.7 = 14
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"11000000000011001100110011001110"), -- -5.8 + 3.6 = -2.2
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000001001011001100110011001101"), -- 9.6 + 1.2 = 10.8
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"01000000001001100110011001100111"), -- 3.9 + -1.3 = 2.6
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111111010011001100110011001100"), -- -2 + 2.8 = 0.8
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"01000000100111001100110011001100"), -- 2.1 + 2.8 = 4.9
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"00111111110011001100110011001100"), -- 7.6 + -6 = 1.6
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"11000001010101001100110011001100"), -- -7.2 + -6.1 = -13.3
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000001001111001100110011001101"), -- -2.2 + -9.6 = -11.8
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000000101100000000000000000000"), -- -2.4 + 7.9 = 5.5
	(b"00111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111111000000000000000000000001"), -- 1.2 + -0.7 = 0.5
	(b"10111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000000100110011001100110011010"), -- -1.3 + 6.1 = 4.8
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000100011001100110011001101"), -- 5.9 + -1.5 = 4.4
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000001000100011001100110011010"), -- -6.3 + -2.8 = -9.1
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000011100110011001100110011"), -- -2.8 + -1 = -3.8
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001010000011001100110011010"), -- -3.6 + -8.5 = -12.1
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001000001001100110011001101"), -- 1.4 + -9.7 = -8.3
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"00111110010011001100110011100000"), -- -7.2 + 7.4 = 0.2
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000001110011001100110011010"), -- 3.2 + -0.3 = 2.9
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"01000000111011001100110011001100"), -- 2.7 + 4.7 = 7.4
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111111001100110011001100110", b"01000000101110011001100110011010"), -- 4 + 1.8 = 5.8
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000001001000000000000000000000"), -- 0.8 + 9.2 = 10
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000000010100110011001100110100"), -- 4.7 + -8 = -3.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000111101100110011001100110"), -- -1 + -6.7 = -7.7
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111111010011001100110011001100"), -- 3.2 + -2.4 = 0.8
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"11000000011011001100110011001100"), -- 0.9 + -4.6 = -3.7
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000000010001100110011001100110"), -- -2.6 + 5.7 = 3.1
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000111111001100110011001100"), -- 8.9 + -1 = 7.9
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"11000000001001100110011001100110"), -- -8.2 + 5.6 = -2.6
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000000010110011001100110011001"), -- 2.3 + -5.7 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101100000000000000000000", b"01000000101100000000000000000000"), -- 0 + 5.5 = 5.5
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000000101011001100110011001101"), -- -0 + 5.4 = 5.4
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"00111110100110011001100110011000"), -- -2.5 + 2.8 = 0.3
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001010110011001100110011001"), -- -9.9 + -3.7 = -13.6
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000111011001100110011001100"), -- 5.1 + 2.3 = 7.4
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"11000000001011001100110011001101"), -- -3.4 + 0.7 = -2.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000001000001100110011001100110"), -- 2.2 + 6.2 = 8.4
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000000100010011001100110011010"), -- 0.6 + -4.9 = -4.3
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"01000000000001100110011001100111"), -- 2.2 + -0.1 = 2.1
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"11000001001001100110011001100110"), -- -9.5 + -0.9 = -10.4
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"10111111000110011001100110011100"), -- 1.8 + -2.4 = -0.6
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001010000011001100110011010"), -- -6.8 + -5.3 = -12.1
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000110000000000000000000000"), -- -1.2 + 7.2 = 6
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000000110111001100110011001101"), -- -0.9 + -6 = -6.9
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000001001010000000000000000000"), -- 4.8 + 5.7 = 10.5
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000001100010100110011001100110"), -- 9.5 + 7.8 = 17.3
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000001000000000000000000000000"), -- -4.5 + -3.5 = -8
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"11000001000011100110011001100111"), -- -1.1 + -7.8 = -8.9
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100011001100110011001101", b"01000000011000000000000000000000"), -- -0.9 + 4.4 = 3.5
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000000111010011001100110011001"), -- -0.9 + 8.2 = 7.3
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000000100100110011001100110100"), -- -3.5 + 8.1 = 4.6
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001011100000000000000000000"), -- 8 + 7 = 15
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000000110010011001100110011010"), -- 0 + 6.3 = 6.3
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"00111111110110011001100110011000"), -- -5.3 + 7 = 1.7
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"01000001011011001100110011001101"), -- 9.8 + 5 = 14.8
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000000110100000000000000000000"), -- -0.1 + -6.4 = -6.5
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000000100100000000000000000000"), -- -4.7 + 9.2 = 4.5
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000000010001100110011001100110"), -- 2.5 + 0.6 = 3.1
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000000100001100110011001100111"), -- -4.4 + 0.2 = -4.2
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"00111111110011001100110011001100"), -- 4.6 + -3 = 1.6
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000111010011001100110011010"), -- -2.5 + -4.8 = -7.3
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000000000011001100110011001100"), -- 7.3 + -9.5 = -2.2
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"01000000100000110011001100110010"), -- 8.9 + -4.8 = 4.1
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"11000000101101100110011001100110"), -- -8.2 + 2.5 = -5.7
	(b"11000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"10111111000110011001100110011000"), -- -7.2 + 6.6 = -0.6
	(b"01000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101001100110011001101", b"11000000111000000000000000000000"), -- 2.3 + -9.3 = -7
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000000010110011001100110011000"), -- 5.5 + -8.9 = -3.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"01000000100010011001100110011010"), -- 0.3 + 4 = 4.3
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000101110011001100110011010"), -- 5 + 0.8 = 5.8
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"11000000101000110011001100110100"), -- -7.4 + 2.3 = -5.1
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000001000111100110011001100110"), -- 9.5 + 0.4 = 9.9
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111001100110011001100110", b"01000000111100110011001100110011"), -- 0.4 + 7.2 = 7.6
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000001000100000000000000000000"), -- 4.4 + 4.6 = 9
	(b"00111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"00111110100110011001100110011010"), -- 1 + -0.7 = 0.3
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000000000001100110011001100100"), -- -6.3 + 8.4 = 2.1
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"00111111011001100110011001100100"), -- -2.7 + 3.6 = 0.9
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111111111001100110011001100110"), -- 2 + -3.8 = -1.8
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"11000001001111100110011001100111"), -- -9.1 + -2.8 = -11.9
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"01000000101101100110011001100111"), -- 0.9 + 4.8 = 5.7
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"11000000001100110011001100110010"), -- -5.2 + 2.4 = -2.8
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000111000000000000000000000"), -- 3.4 + 3.6 = 7
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"01000000100101100110011001100111"), -- -3.6 + 8.3 = 4.7
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001100000110011001100110011"), -- 9.4 + 7 = 16.4
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001100001110011001100110011"), -- -9.3 + -7.6 = -16.9
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"10111111010011001100110011010000"), -- 8.7 + -9.5 = -0.8
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000001010110000000000000000000"), -- -9.1 + -4.4 = -13.5
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000000101100110011001100110100"), -- 4 + -9.6 = -5.6
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000001001010000000000000000000"), -- -3.2 + -7.3 = -10.5
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100010011001100110011010", b"10111111110000000000000000000000"), -- -5.8 + 4.3 = -1.5
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"11000000001111111111111111111110"), -- 5.9 + -8.9 = -3
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000000001000000000000000000000"), -- -4.5 + 7 = 2.5
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"11000000000110011001100110011000"), -- -7.7 + 5.3 = -2.4
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000100000000000000000000", b"01000001000101001100110011001101"), -- 0.3 + 9 = 9.3
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000000100110011001100110011010"), -- 4.7 + -9.5 = -4.8
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"11000001001010000000000000000000"), -- -3.4 + -7.1 = -10.5
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"01000000111010011001100110011010"), -- 8.3 + -1 = 7.3
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"01000000000000000000000000000000"), -- 6.4 + -4.4 = 2
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"01000000011001100110011001100110"), -- 7.7 + -4.1 = 3.6
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"10111110100110011001100110010000"), -- -8.2 + 7.9 = -0.3
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"00111111111100110011001100110100"), -- 7.5 + -5.6 = 1.9
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000001001110000000000000000000"), -- 8.8 + 2.7 = 11.5
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000000101000000000000000000000"), -- 4.8 + -9.8 = -5
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"01000000111011001100110011001100"), -- 2.7 + 4.7 = 7.4
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"01000000100100000000000000000001"), -- -4.1 + 8.6 = 4.5
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"10111111110000000000000000000000"), -- 4.6 + -6.1 = -1.5
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000000000011001100110011001100"), -- 7.3 + -9.5 = -2.2
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000000001001100110011001101000"), -- -5.2 + 7.8 = 2.6
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"10111111001100110011001100111000"), -- -6.3 + 5.6 = -0.7
	(b"00111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000000111011001100110011001101"), -- 1.1 + 6.3 = 7.4
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000000000000000000000000000000"), -- 6.5 + -8.5 = -2
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111111110110011001100110011010"), -- -2.5 + 0.8 = -1.7
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"00111111110110011001100110011100"), -- 4.8 + -3.1 = 1.7
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001010111100110011001100110"), -- -7.6 + -6.3 = -13.9
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001001011100110011001100110"), -- -5.2 + -5.7 = -10.9
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000001010110110011001100110100"), -- 5.9 + 7.8 = 13.7
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000001001110011001100110011001"), -- 8.4 + 3.2 = 11.6
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001011110011001100110011010"), -- -7.6 + -8 = -15.6
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"10111110010011001100110011000000"), -- 9.2 + -9.4 = -0.2
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000001000010011001100110011010"), -- -6.8 + -1.8 = -8.6
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000011000000000000000000000"), -- -2.5 + -1 = -3.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"10111111010011001100110011001110"), -- 0.4 + -1.2 = -0.8
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000001000011100110011001100110"), -- -7.1 + -1.8 = -8.9
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"01000000011110011001100110011100"), -- 8.1 + -4.2 = 3.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101100000000000000000000", b"01000000101001100110011001100110"), -- -0.3 + 5.5 = 5.2
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000000001111111111111111111110"), -- -5.4 + 8.4 = 3
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"01000001000000000000000000000000"), -- 4 + 4 = 8
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"11000000010100110011001100110100"), -- -8.6 + 5.3 = -3.3
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000011100110011001100110011"), -- 0.1 + 3.7 = 3.8
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000001011011100110011001100110"), -- -7.7 + -7.2 = -14.9
	(b"01000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"10111111100000000000000000000000"), -- 4.1 + -5.1 = -1
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000110001100110011001100111"), -- 0.6 + -6.8 = -6.2
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000001011010000000000000000000"), -- -7.9 + -6.6 = -14.5
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000001001101100110011001100110"), -- -7.3 + -4.1 = -11.4
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001011011001100110011001100"), -- 8.7 + 6.1 = 14.8
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000001011111100110011001100110"), -- -8.7 + -7.2 = -15.9
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"11000000110001100110011001100110"), -- -6.2 + -0 = -6.2
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000000010011001100110011001100"), -- -6.7 + 9.9 = 3.2
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"10111111111001100110011001101000"), -- -6.3 + 4.5 = -1.8
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000000100010011001100110011001"), -- 5.1 + -9.4 = -4.3
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"10111111100000000000000000000000"), -- 0.7 + -1.7 = -1
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"10111111100110011001100110011010"), -- -5 + 3.8 = -1.2
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"10111111111001100110011001100110"), -- -3.1 + 1.3 = -1.8
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000000000000000000000000000"), -- -2.5 + 0.5 = -2
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000001000001001100110011001100"), -- -1.1 + 9.4 = 8.3
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000001000000110011001100110011"), -- 7.2 + 1 = 8.2
	(b"11000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"11000000000110011001100110011010"), -- -7.4 + 5 = -2.4
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"00111111110011001100110011010000"), -- 9.8 + -8.2 = 1.6
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"11000000001001100110011001100110"), -- -9 + 6.4 = -2.6
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"00111111100011001100110011001000"), -- 9.2 + -8.1 = 1.1
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"10111111011001100110011001101000"), -- 5.6 + -6.5 = -0.9
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000001011010000000000000000000"), -- 4.6 + 9.9 = 14.5
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000000011000000000000000000000"), -- -1.9 + 5.4 = 3.5
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"11000000110111001100110011001101"), -- -2.1 + -4.8 = -6.9
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000000111010011001100110011010"), -- 1.5 + -8.8 = -7.3
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000000110110011001100110011010"), -- 4.9 + 1.9 = 6.8
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"00111111000110011001100110011000"), -- 5.1 + -4.5 = 0.6
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"10111111101001100110011001100111"), -- 0.9 + -2.2 = -1.3
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000001000101001100110011001101"), -- 9.6 + -0.3 = 9.3
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000001100110011001100110", b"01000001001011001100110011001100"), -- 2.4 + 8.4 = 10.8
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000001010110110011001100110100"), -- -5.6 + -8.1 = -13.7
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"01000000110101100110011001100110"), -- 9.2 + -2.5 = 6.7
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"00111111101001100110011001101000"), -- -8.3 + 9.6 = 1.3
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"01000000111001100110011001100110"), -- -0.8 + 8 = 7.2
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001001011100110011001100110"), -- -5.6 + -5.3 = -10.9
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000000100111001100110011001101"), -- -2 + -2.9 = -4.9
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"), -- 6.3 + -6.3 = 0
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"01000001011110000000000000000000"), -- 6.9 + 8.6 = 15.5
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"01000001000010011001100110011010"), -- 5.5 + 3.1 = 8.6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000010000000000000000000000"), -- 0.8 + -3.8 = -3
	(b"11000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001010010000000000000000000"), -- -6.8 + -5.7 = -12.5
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"01000000101110011001100110011010"), -- -2.2 + 8 = 5.8
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100011001100110011001101", b"01000001000001100110011001100110"), -- 4 + 4.4 = 8.4
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000001010011100110011001100111"), -- 9.6 + 3.3 = 12.9
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001001100011001100110011010"), -- -2.9 + -8.2 = -11.1
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"10111111101001100110011001100111"), -- 1.9 + -3.2 = -1.3
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000001001010110011001100110011"), -- 7 + 3.7 = 10.7
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010000000000000000000000", b"11000000100100000000000000000000"), -- -1.5 + -3 = -4.5
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"01000000101000110011001100110011"), -- 5.6 + -0.5 = 5.1
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000001110011001100110011010"), -- -1.9 + -1 = -2.9
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000001010111100110011001100110"), -- -7.9 + -6 = -13.9
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000000010100110011001100110011"), -- -3.2 + 6.5 = 3.3
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"00111101110011001100110011000000"), -- 2.5 + -2.4 = 0.0999999
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"01000000100001100110011001100111"), -- 8.8 + -4.6 = 4.2
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000000010000000000000000000000"), -- -2.3 + -0.7 = -3
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"01000000001011001100110011001110"), -- -4.2 + 6.9 = 2.7
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000001011000011001100110011010"), -- 6.2 + 7.9 = 14.1
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"01000000010001100110011001101000"), -- 8.8 + -5.7 = 3.1
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000000101010011001100110011010"), -- 2.7 + -8 = -5.3
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"01000000100011001100110011001100"), -- -2.3 + 6.7 = 4.4
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000111100110011001100110", b"11000000010110011001100110011000"), -- 6.5 + -9.9 = -3.4
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000001100001000000000000000000"), -- 7.6 + 8.9 = 16.5
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000010110011001100110011001"), -- -0.8 + 4.2 = 3.4
	(b"01000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000111100110011001100110011"), -- 6.6 + 1 = 7.6
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000001011000110011001100110011"), -- 8 + 6.2 = 14.2
	(b"11000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"00111111000000000000000000000000"), -- -7.3 + 7.8 = 0.5
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000001011011100110011001100110"), -- 8.4 + 6.5 = 14.9
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000111011001100110011001101"), -- -4.9 + -2.5 = -7.4
	(b"01000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"01000000011100110011001100110011"), -- 5 + -1.2 = 3.8
	(b"11000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000001001010000000000000000000"), -- -5.2 + -5.3 = -10.5
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"11000000010110011001100110011010"), -- -7 + 3.6 = -3.4
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000000100000110011001100110011"), -- 1.4 + 2.7 = 4.1
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000001000100110011001100110011"), -- 3.5 + 5.7 = 9.2
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"11000001010100011001100110011010"), -- -8.5 + -4.6 = -13.1
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000000100100000000000000000000"), -- -5.7 + 1.2 = -4.5
	(b"11000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001001100011001100110011010"), -- -4.8 + -6.3 = -11.1
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010001100110011001100110", b"11000000000110011001100110011010"), -- -5.5 + 3.1 = -2.4
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000000110000110011001100110010"), -- 3.3 + -9.4 = -6.1
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000001000001100110011001100110"), -- -9.7 + 1.3 = -8.4
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001010011100110011001100110"), -- -9.2 + -3.7 = -12.9
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000000101001100110011001100111"), -- 4.3 + 0.9 = 5.2
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000001000100011001100110011010"), -- -0.1 + -9 = -9.1
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000000100101100110011001100110"), -- -2.7 + 7.4 = 4.7
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001011001100110011001101", b"01000000001100110011001100110011"), -- 5.5 + -2.7 = 2.8
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"01000000001011001100110011001100"), -- 4.2 + -1.5 = 2.7
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"01000000001110011001100110011010"), -- 1.3 + 1.6 = 2.9
	(b"11000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"00111101110011001100110010000000"), -- -8.1 + 8.2 = 0.0999994
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"00111110110011001100110011001000"), -- 3.8 + -3.4 = 0.4
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"00111111110110011001100110011010"), -- 0.7 + 1 = 1.7
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000100100000000000000000000"), -- 3 + 1.5 = 4.5
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"11000000110111001100110011001110"), -- -8.6 + 1.7 = -6.9
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000001010011001100110011001100"), -- 3.6 + 9.2 = 12.8
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"01000000111111001100110011001101"), -- 2.6 + 5.3 = 7.9
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"11000000000011001100110011001100"), -- -4.1 + 1.9 = -2.2
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001000101100110011001100110"), -- -0.7 + -8.7 = -9.4
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000000011100110011001100110011"), -- 1.5 + 2.3 = 3.8
	(b"01000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"10111111100110011001100110011000"), -- 7.7 + -8.9 = -1.2
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"11000001000011100110011001100110"), -- -2.9 + -6 = -8.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000001000100110011001100110011"), -- 3 + 6.2 = 9.2
	(b"00111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001000101100110011001100110"), -- 0.3 + -9.7 = -9.4
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000001000111001100110011001101"), -- 9.1 + 0.7 = 9.8
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000000101101100110011001100111"), -- 0.1 + -5.8 = -5.7
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"10111111110000000000000000000000"), -- -8.2 + 6.7 = -1.5
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000001001001100110011001100110"), -- -4 + -6.4 = -10.4
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"11000001001010011001100110011010"), -- -6.6 + -4 = -10.6
	(b"01000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000001001000011001100110011010"), -- 8.6 + 1.5 = 10.1
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000000010011001100110011001110"), -- -5.9 + 9.1 = 3.2
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000000000001100110011001100110"), -- -2.1 + 4.2 = 2.1
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"01000001001110110011001100110011"), -- 7.5 + 4.2 = 11.7
	(b"10111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"00111110010011001100110011010000"), -- -1.8 + 2 = 0.2
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000110110011001100110011001"), -- 4.7 + 2.1 = 6.8
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000001100001110011001100110100"), -- -9.6 + -7.3 = -16.9
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"01000001001110110011001100110011"), -- 7.1 + 4.6 = 11.7
	(b"10111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000001000001100110011001100111"), -- -0.7 + 9.1 = 8.4
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110011001100110011001101", b"00111111100110011001100110011010"), -- -0.4 + 1.6 = 1.2
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000000110010011001100110011010"), -- 1.8 + -8.1 = -6.3
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000011001100110011001100110"), -- -2 + -1.6 = -3.6
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"00111110110011001100110011010000"), -- 2.2 + -1.8 = 0.4
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000001100001011001100110011010"), -- 6.8 + 9.9 = 16.7
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"11000000101001100110011001100110"), -- -2.7 + -2.5 = -5.2
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000001000111001100110011001101"), -- -9.6 + -0.2 = -9.8
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"00111101110011001100110011000000"), -- 7.1 + -7 = 0.0999999
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000000101001100110011001100110"), -- -3.1 + -2.1 = -5.2
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000001000100011001100110011010"), -- -0.6 + -8.5 = -9.1
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"10111111000000000000000000000000"), -- -7.1 + 6.6 = -0.5
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000000010000000000000000000000"), -- -3.6 + 0.6 = -3
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000110011001100110011010", b"11000000110001100110011001100111"), -- -8.6 + 2.4 = -6.2
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001000000110011001100110011"), -- -3.7 + -4.5 = -8.2
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"00111111110011001100110011001100"), -- -5.1 + 6.7 = 1.6
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"11000000011011001100110011001101"), -- -2.7 + -1 = -3.7
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000001001010011001100110011010"), -- -1 + -9.6 = -10.6
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"), -- -1.5 + 1.5 = 0
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100000110011001100110011", b"01000000011001100110011001100110"), -- -0.5 + 4.1 = 3.6
	(b"00111111101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"01000001000110011001100110011010"), -- 1.3 + 8.3 = 9.6
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000000101101100110011001100110"), -- -4.2 + -1.5 = -5.7
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"10111110110011001100110011010000"), -- -3.2 + 2.8 = -0.4
	(b"11000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000000111000000000000000000000"), -- -2.2 + 9.2 = 7
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100101100110011001100110", b"11000000010000000000000000000000"), -- -7.7 + 4.7 = -3
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"00111111000000000000000000000000"), -- 9.5 + -9 = 0.5
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001010011100110011001100110"), -- -7.7 + -5.2 = -12.9
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"11000000001001100110011001101000"), -- -9.3 + 6.7 = -2.6
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"11000001001010110011001100110100"), -- -8.6 + -2.1 = -10.7
	(b"01000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000000001110011001100110011001"), -- 3.3 + -6.2 = -2.9
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000001000000110011001100110011"), -- -1.2 + 9.4 = 8.2
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"01000000101011001100110011001100"), -- -3.8 + 9.2 = 5.4
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"11000001000111001100110011001101"), -- -3.5 + -6.3 = -9.8
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100011001100110011010", b"01000001000101001100110011001101"), -- 0.2 + 9.1 = 9.3
	(b"01000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"11000000011110011001100110011100"), -- 4.2 + -8.1 = -3.9
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000000110110011001100110011001"), -- 2.4 + -9.2 = -6.8
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"11000000111101100110011001100110"), -- -6.6 + -1.1 = -7.7
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000000000001100110011001100110"), -- 1.6 + -3.7 = -2.1
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111100000000000000000000000", b"01000000110000110011001100110011"), -- 5.1 + 1 = 6.1
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"01000000110010011001100110011001"), -- 8.4 + -2.1 = 6.3
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001100000011001100110011010"), -- -8.3 + -7.9 = -16.2
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"00111110110011001100110011010000"), -- -5.9 + 6.3 = 0.4
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000001001100000000000000000000"), -- 9.8 + 1.2 = 11
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000000111111001100110011001101"), -- 0.6 + 7.3 = 7.9
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000001000010000000000000000000"), -- 5.3 + 3.2 = 8.5
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100101100110011001100110", b"11000001000100000000000000000000"), -- -4.3 + -4.7 = -9
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"11000000000100110011001100110100"), -- -7.9 + 5.6 = -2.3
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000001010000110011001100110100"), -- -2.4 + -9.8 = -12.2
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"01000000110010011001100110011010"), -- 8.3 + -2 = 6.3
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"11000000001011001100110011001110"), -- -8.6 + 5.9 = -2.7
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000000110110011001100110011001"), -- 7.1 + -0.3 = 6.8
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000001001010000000000000000000"), -- -9.3 + -1.2 = -10.5
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000001000000000000000000000000"), -- -4.9 + -3.1 = -8
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000000101110011001100110011010"), -- 3.6 + 2.2 = 5.8
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000001001100110011001100110"), -- 2.8 + -0.2 = 2.6
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000001010010110011001100110100"), -- -9.6 + -3.1 = -12.7
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"11000001001000110011001100110011"), -- -0.5 + -9.7 = -10.2
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000000110000110011001100110100"), -- -2.7 + 8.8 = 6.1
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"10111111110000000000000000000000"), -- 4.4 + -5.9 = -1.5
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110000110011001100110011", b"11000000110011001100110011001101"), -- -0.3 + -6.1 = -6.4
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000000110101100110011001100110"), -- 3 + 3.7 = 6.7
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"11000000001110011001100110011001"), -- 0.2 + -3.1 = -2.9
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"00111111000000000000000000000000"), -- -6 + 6.5 = 0.5
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"01000001000000000000000000000000"), -- 5.4 + 2.6 = 8
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"10111111011001100110011001100000"), -- -9.5 + 8.6 = -0.9
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000001010100011001100110011001"), -- -9.4 + -3.7 = -13.1
	(b"11000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"00111111110110011001100110011000"), -- -4.8 + 6.5 = 1.7
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001000100000000000000000000"), -- -3.3 + -5.7 = -9
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000000101110011001100110011001"), -- -0.6 + -5.2 = -5.8
	(b"10111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000000101011001100110011001100"), -- -0.8 + 6.2 = 5.4
	(b"11000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001001001100110011001100110"), -- -2.5 + -7.9 = -10.4
	(b"01000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000101010011001100110011001"), -- 5.2 + 0.1 = 5.3
	(b"10111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"01000001000011100110011001100110"), -- -0.6 + 9.5 = 8.9
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101000110011001100110011", b"01000001000110000000000000000000"), -- 4.4 + 5.1 = 9.5
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"01000000100100110011001100110011"), -- 8.7 + -4.1 = 4.6
	(b"11000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"11000001010111001100110011001100"), -- -7.6 + -6.2 = -13.8
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000000000011001100110011001100"), -- 7.2 + -9.4 = -2.2
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111000110011001100110011010", b"11000000101000000000000000000000"), -- -4.4 + -0.6 = -5
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000001001000110011001100110011"), -- 1.4 + 8.8 = 10.2
	(b"01000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001011000011001100110011010"), -- 8 + 6.1 = 14.1
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"00111111100110011001100110011010"), -- -2.8 + 4 = 1.2
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000111100110011001100110011"), -- -0.9 + -6.7 = -7.6
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110000110011001100110011", b"01000001011000110011001100110100"), -- 8.1 + 6.1 = 14.2
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"01000001001011100110011001100110"), -- 2.9 + 8 = 10.9
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"10111111110011001100110011001000"), -- -9.4 + 7.8 = -1.6
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000000110110011001100110011010"), -- -1 + -5.8 = -6.8
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000000101000110011001100110011"), -- -4.6 + 9.7 = 5.1
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"11000000000110011001100110011010"), -- -7.8 + 5.4 = -2.4
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"01000000010100110011001100110100"), -- 9.6 + -6.3 = 3.3
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"10111111011001100110011001101000"), -- 3.9 + -4.8 = -0.9
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000000110110011001100110011010"), -- 4.3 + 2.5 = 6.8
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000001001100110011001100110100"), -- -3.9 + -7.3 = -11.2
	(b"01000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110011001100110011001101", b"01000001011010110011001100110100"), -- 8.3 + 6.4 = 14.7
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000000000110011001100110011001"), -- 1.7 + -4.1 = -2.4
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"01000000101000110011001100110010"), -- 8.4 + -3.3 = 5.1
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000001000001001100110011001101"), -- -9.7 + 1.4 = -8.3
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000010000000000000000000001"), -- 3.8 + -6.8 = -3
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000000011001100110011001100110"), -- 4 + -0.4 = 3.6
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"01000000010001100110011001100110"), -- -1.4 + 4.5 = 3.1
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"01000000110011001100110011001101"), -- 6.3 + 0.1 = 6.4
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000001001111100110011001100110"), -- -8.3 + -3.6 = -11.9
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000011110011001100110011010"), -- 2.9 + -6.8 = -3.9
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000001000110000000000000000000"), -- -1.1 + -8.4 = -9.5
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000000000011001100110011001100"), -- -1.4 + 3.6 = 2.2
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000000101000110011001100110100"), -- 2.2 + -7.3 = -5.1
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000000100101100110011001100111"), -- -1.1 + 5.8 = 4.7
	(b"11000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001000001001100110011001100"), -- -3.1 + -5.2 = -8.3
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000001100110011001100110", b"00111110100110011001100110100000"), -- 2.4 + -2.1 = 0.3
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000100110011001100110011", b"00111111011001100110011001100000"), -- -8.3 + 9.2 = 0.9
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010001100110011001100110", b"00111111100110011001100110011100"), -- 4.3 + -3.1 = 1.2
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000000101111001100110011001101"), -- 2.4 + -8.3 = -5.9
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001001011100110011001100110"), -- -5.7 + -5.2 = -10.9
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111011001100110011001100110", b"01000000111100110011001100110011"), -- 8.5 + -0.9 = 7.6
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111110000000000000000000000", b"01000000100100000000000000000000"), -- 3 + 1.5 = 4.5
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000000101001100110011001100110"), -- -2.6 + -2.6 = -5.2
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"01000000000110011001100110011010"), -- -3.9 + 6.3 = 2.4
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101000000000000000000000", b"10111111110110011001100110011000"), -- -6.7 + 5 = -1.7
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"01000001010011100110011001100110"), -- 6.4 + 6.5 = 12.9
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"01000000101001100110011001100110"), -- 8.4 + -3.2 = 5.2
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"01000000010000000000000000000000"), -- 5.6 + -2.6 = 3
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000000000000000000000", b"10111111100000000000000000000000"), -- -9 + 8 = -1
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111100110011001100110011", b"01000000110000110011001100110011"), -- -1.5 + 7.6 = 6.1
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110001100110011001100110", b"00111111111100110011001100111000"), -- 8.1 + -6.2 = 1.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000000110001100110011001100110"), -- 2.8 + -9 = -6.2
	(b"01000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000001001010000000000000000000"), -- 7.1 + 3.4 = 10.5
	(b"00111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000000111110011001100110011010"), -- 0.2 + -8 = -7.8
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"11000001000100000000000000000000"), -- 0.1 + -9.1 = -9
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000001010000011001100110011010"), -- -3.9 + -8.2 = -12.1
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000001000000000000000000000", b"01000001000001100110011001100110"), -- 5.9 + 2.5 = 8.4
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000000000000000000000000", b"00111111110011001100110011001100"), -- 3.6 + -2 = 1.6
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"01000001011001001100110011001101"), -- 9.5 + 4.8 = 14.3
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000100010011001100110011010", b"10111111010011001100110011001000"), -- -5.1 + 4.3 = -0.8
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000001010110110011001100110011"), -- -7.1 + -6.6 = -13.7
	(b"11000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000000000110011001100110011010"), -- -2.9 + 0.5 = -2.4
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001001110011001100110011010"), -- -3.6 + -8 = -11.6
	(b"00111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000001000101100110011001100111"), -- 1.6 + 7.8 = 9.4
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"10111111110110011001100110011010"), -- 1.8 + -3.5 = -1.7
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000000010011001100110011001101"), -- 2.2 + -5.4 = -3.2
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"11000000000001100110011001100110"), -- -8 + 5.9 = -2.1
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000001000000110011001100110011"), -- 6.2 + 2 = 8.2
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"00111111100000000000000000000000"), -- 5.8 + -4.8 = 1
	(b"01000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"10111101110011001100110011000000"), -- 5.5 + -5.6 = -0.0999999
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101101100110011001100110", b"11000001000100011001100110011010"), -- -3.4 + -5.7 = -9.1
	(b"11000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000000111111001100110011001101"), -- -2.6 + -5.3 = -7.9
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000000011100110011001100110100"), -- 0.4 + 3.4 = 3.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000000101110011001100110011010"), -- -0 + -5.8 = -5.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000000100100000000000000000000"), -- 3.8 + 0.7 = 4.5
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000001001110110011001100110011"), -- 9.8 + 1.9 = 11.7
	(b"00111111001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001000011001100110011001101"), -- 0.7 + -9.5 = -8.8
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"11000000010001100110011001100111"), -- 3.8 + -6.9 = -3.1
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000110110011001100110011", b"01000000100100110011001100110011"), -- -5.1 + 9.7 = 4.6
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000010011001100110011010", b"01000001100011100110011001100110"), -- 9.2 + 8.6 = 17.8
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"11000000110110011001100110011001"), -- -6.6 + -0.2 = -6.8
	(b"00111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000000111000000000000000000000"), -- 1.7 + -8.7 = -7
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"01000000010100110011001100110100"), -- 7.5 + -4.2 = 3.3
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000001011011100110011001100110"), -- 7.6 + 7.3 = 14.9
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000011001100110011001101", b"11000001100010100110011001100110"), -- -8.5 + -8.8 = -17.3
	(b"01000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000000001110011001100110011000"), -- 4.3 + -7.2 = -2.9
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000000010011001100110011001101"), -- -0 + 3.2 = 3.2
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"10111110010011001100110100000000"), -- 8.9 + -9.1 = -0.200001
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"01000000110000110011001100110011"), -- 2.6 + 3.5 = 6.1
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000110010011001100110011010"), -- -4.9 + -1.4 = -6.3
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000001010001001100110011001100"), -- -4.7 + -7.6 = -12.3
	(b"01000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110000000000000000000000", b"01000000000110011001100110011000"), -- 8.4 + -6 = 2.4
	(b"11000000111101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100100000000000000000000", b"11000001010000110011001100110011"), -- -7.7 + -4.5 = -12.2
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"11000000100000110011001100110100"), -- 2.7 + -6.8 = -4.1
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010110011001100110011010", b"01000001001111100110011001100110"), -- 8.5 + 3.4 = 11.9
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000000101000000000000000000000"), -- -1.5 + -3.5 = -5
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111010011001100110011010", b"11000001011111001100110011001101"), -- -8.5 + -7.3 = -15.8
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000111001100110011001100110"), -- -6 + -1.2 = -7.2
	(b"11000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"11000000101110011001100110011010"), -- -9.1 + 3.3 = -5.8
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"01000000001110011001100110011010"), -- 8.5 + -5.6 = 2.9
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000000101000110011001100110100"), -- -2.3 + 7.4 = 5.1
	(b"01000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"11000000100011001100110011001100"), -- 2.7 + -7.1 = -4.4
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"00111111100011001100110011001100"), -- 6.9 + -5.8 = 1.1
	(b"01000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"01000000000001100110011001100110"), -- 9 + -6.9 = 2.1
	(b"01000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"01000000001011001100110011001101"), -- 6 + -3.3 = 2.7
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000001011011100110011001100110"), -- -8.5 + -6.4 = -14.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100110011001100110011010", b"10111111111001100110011001101000"), -- 3 + -4.8 = -1.8
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"11000000010110011001100110011001"), -- 2.2 + -5.6 = -3.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"01000000110000000000000000000000"), -- 0 + 6 = 6
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"10111101110011001100110011001000"), -- -0.9 + 0.8 = -0.1
	(b"01000000001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"11000000001001100110011001100110"), -- 2.9 + -5.5 = -2.6
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"11000000110111001100110011001101"), -- -5 + -1.9 = -6.9
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000000101111001100110011001101"), -- -3.5 + -2.4 = -5.9
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000001000011100110011001100110"), -- -6.6 + -2.3 = -8.9
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"11000000111001100110011001100110"), -- -5.6 + -1.6 = -7.2
	(b"11000000001011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"11000001000000110011001100110011"), -- -2.7 + -5.5 = -8.2
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101100000000000000000000", b"01000000100001100110011001100110"), -- 9.7 + -5.5 = 4.2
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"), -- 1.5 + -1.5 = 0
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"01000000010100110011001100110100"), -- -1.6 + 4.9 = 3.3
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000001001100000000000000000000"), -- -4.6 + -6.4 = -11
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"01000000110000110011001100110011"), -- 5.9 + 0.2 = 6.1
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"01000000100010011001100110011010"), -- 6.1 + -1.8 = 4.3
	(b"01000000010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"00111111010011001100110011001100"), -- 3.1 + -2.3 = 0.8
	(b"01000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"01000000000001100110011001100110"), -- 4.5 + -2.4 = 2.1
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000001010011001100110011001101"), -- 7 + 5.8 = 12.8
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"01000000000011001100110011001100"), -- 0.1 + 2.1 = 2.2
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000000001110011001100110011010"), -- -3.9 + 6.8 = 2.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111100000000000000000000000", b"00111111111001100110011001100110"), -- 2.8 + -1 = 1.8
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"00111111111100110011001100111000"), -- 9.1 + -7.2 = 1.9
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111011001100110011001101", b"01000001010110000000000000000000"), -- 6.1 + 7.4 = 13.5
	(b"01000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"01000000101000110011001100110010"), -- 8.9 + -3.8 = 5.1
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"01000000110111001100110011001100"), -- 8.7 + -1.8 = 6.9
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"11000001010001001100110011001100"), -- -7.1 + -5.2 = -12.3
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"11000001001010000000000000000000"), -- -6.4 + -4.1 = -10.5
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000001001001100110011001100110"), -- -6.6 + -3.8 = -10.4
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"01000000100011001100110011001110"), -- 9.6 + -5.2 = 4.4
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000000000000000000000000", b"11000001011011100110011001100110"), -- -6.9 + -8 = -14.9
	(b"01000000111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101000000000000000000000", b"01000000000100110011001100110100"), -- 7.3 + -5 = 2.3
	(b"11000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101011001100110011001101", b"01000000001001100110011001100111"), -- -2.8 + 5.4 = 2.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000000010100110011001100110011"), -- 3.5 + -0.2 = 3.3
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110011001100110011001101", b"11000000001000000000000000000000"), -- 3.9 + -6.4 = -2.5
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"01000001100000110011001100110011"), -- 9.4 + 7 = 16.4
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111110110011001100110011001000"), -- 3.4 + -3.8 = -0.4
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"00111111010011001100110011001000"), -- -5.8 + 6.6 = 0.8
	(b"01000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000001100110011001100110", b"11000000000111111111111111111110"), -- 5.9 + -8.4 = -2.5
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"10111111000110011001100110011100"), -- 2.8 + -3.4 = -0.6
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000001001111001100110011001101"), -- -9.6 + -2.2 = -11.8
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000000110000110011001100110011"), -- 4.7 + 1.4 = 6.1
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"10111111001100110011001100110100"), -- 2.6 + -3.3 = -0.7
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"01000000101001100110011001100111"), -- 4.4 + 0.8 = 5.2
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"01000000001011001100110011001100"), -- -3.9 + 6.6 = 2.7
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"10111111010011001100110011010000"), -- 8.7 + -9.5 = -0.8
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"10111111101001100110011001101000"), -- 3 + -4.3 = -1.3
	(b"01000001000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000001001011001100110011001101"), -- 8.1 + 2.7 = 10.8
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000000110110011001100110011010"), -- -5.4 + -1.4 = -6.8
	(b"01000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"01000000011110011001100110011010"), -- 8.8 + -4.9 = 3.9
	(b"01000000111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000001010101100110011001100110"), -- 7.6 + 5.8 = 13.4
	(b"11000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000101010011001100110011010", b"10111111100011001100110011001100"), -- -6.4 + 5.3 = -1.1
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011100110011001100110011", b"00111110110011001100110011001000"), -- -3.4 + 3.8 = 0.4
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"), -- 4 + -4 = 0
	(b"01000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"10111110010011001100110011010000"), -- 3.6 + -3.8 = -0.2
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"11000000000001100110011001101000"), -- 7.5 + -9.6 = -2.1
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010110011001100110011", b"11000001100011001100110011001100"), -- -8.9 + -8.7 = -17.6
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000001010101001100110011001100"), -- 4.4 + 8.9 = 13.3
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000001000000110011001100110011"), -- -3.8 + -4.4 = -8.2
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000011000000000000000000000", b"11000000101000000000000000000000"), -- -8.5 + 3.5 = -5
	(b"01000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000001011101001100110011001100"), -- 9.7 + 5.6 = 15.3
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"01000000001100110011001100110011"), -- -0.2 + 3 = 2.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000000011110011001100110011001"), -- 3.7 + -7.6 = -3.9
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100011001100110011001101", b"11000000100100110011001100110011"), -- -9 + 4.4 = -4.6
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000001000111001100110011001101"), -- 1.9 + 7.9 = 9.8
	(b"01000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000001010010000000000000000000"), -- 3.7 + 8.8 = 12.5
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"11000001000000000000000000000000"), -- -4 + -4 = -8
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"10111101110011001100110011001110"), -- -0.3 + 0.2 = -0.1
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100100110011001100110011", b"11000000100000000000000000000001"), -- -8.6 + 4.6 = -4
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111011001100110011001101", b"11000001010111100110011001100110"), -- -6.5 + -7.4 = -13.9
	(b"11000001000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000001001111100110011001100110"), -- -8 + -3.9 = -11.9
	(b"01000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000000100110011001100110011010"), -- 4.4 + 0.4 = 4.8
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000111101100110011001100110", b"11000001001110110011001100110011"), -- -4 + -7.7 = -11.7
	(b"01000001000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"01000000000000000000000000000010"), -- 9.1 + -7.1 = 2
	(b"00111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011110011001100110011010", b"01000000101010011001100110011010"), -- 1.4 + 3.9 = 5.3
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000001000001001100110011001101"), -- 7.8 + 0.5 = 8.3
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"01000001000010110011001100110011"), -- 7.8 + 0.9 = 8.7
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"00111110010011001100110011000000"), -- -4 + 4.2 = 0.2
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"11000001100101011001100110011010"), -- -9.3 + -9.4 = -18.7
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"11000000010011001100110011001100"), -- -0.9 + -2.3 = -3.2
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000010011001100110011001101", b"11000001001110110011001100110011"), -- -8.5 + -3.2 = -11.7
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"11000001000001100110011001100110"), -- 0.8 + -9.2 = -8.4
	(b"01000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"01000001000110000000000000000000"), -- 3.9 + 5.6 = 9.5
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"01000000011000000000000000000000"), -- -4.4 + 7.9 = 3.5

	(b"11000010001101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001100011001100110011010", b"10111111100110011001100110000000"), -- -45.6 + 44.4 = -1.2
	(b"11000010001010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110010011001100110011010", b"11000010000011111001100110011010"), -- -42.2 + 6.3 = -35.9
	(b"01000001110101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000100010011001100110011", b"01000010011110111001100110011010"), -- 26.6 + 36.3 = 62.9
	(b"01000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"01000001001100110011001100110011"), -- 9.2 + 2 = 11.2
	(b"11000010110000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001100000000000000000", b"11000001010111001100110011010000"), -- -96.8 + 83 = -13.8
	(b"11000010100111101001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100100111100110011001101", b"11000011000110010011001100110100"), -- -79.3 + -73.9 = -153.2
	(b"11000010100001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010100100110011001100110", b"11000010111011010011001100110011"), -- -66 + -52.6 = -118.6
	(b"11000010101001100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010000110011001100110", b"11000001011011100110011001101000"), -- -83.1 + 68.2 = -14.9
	(b"11000010001101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001110011001100110011010", b"11000010101101111100110011001101"), -- -45.5 + -46.4 = -91.9
	(b"01000010100001110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001000010011001100110011", b"01000001110110110011001100110010"), -- 67.7 + -40.3 = 27.4
	(b"11000010011011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011101011001100110011010", b"00111111110011001100110011100000"), -- -59.8 + 61.4 = 1.6
	(b"11000010000110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100111100110011001101", b"11000010111000000110011001100110"), -- -38.3 + -73.9 = -112.2
	(b"11000010100101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111011011001100110011010", b"11000010001100101100110011001101"), -- -74.4 + 29.7 = -44.7
	(b"01000001111100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100010100011001100110011", b"11000010000110110011001100110011"), -- 30.3 + -69.1 = -38.8
	(b"01000010100111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011010000110011001100110", b"01000011000010011011001100110011"), -- 79.6 + 58.1 = 137.7
	(b"11000001101001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000011111001100110011010", b"01000001011100000000000000000010"), -- -20.9 + 35.9 = 15
	(b"01000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101110000000000000000", b"11000010101100000011001100110011"), -- 3.4 + -91.5 = -88.1
	(b"11000010000100010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000110100110011001100110", b"11000010100101011100110011001100"), -- -36.3 + -38.6 = -74.9
	(b"01000010000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100001100110011001101", b"11000010000001100110011001100111"), -- 38.8 + -72.4 = -33.6
	(b"01000001001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100001011001100110011010", b"01000010100110111100110011001101"), -- 11.1 + 66.8 = 77.9
	(b"01000010001011010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101000110000000000000000", b"11000010000110001100110011001101"), -- 43.3 + -81.5 = -38.2
	(b"11000010110001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010100000000000000000", b"11000001111011001100110011001100"), -- -98.6 + 69 = -29.6
	(b"11000010001000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100000101001100110011010", b"11000010110100101100110011001101"), -- -40.1 + -65.3 = -105.4
	(b"01000010011011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101010101100110011001101", b"01000011000100010001100110011010"), -- 59.7 + 85.4 = 145.1
	(b"01000010001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110001100110011001101", b"01000010111011000000000000000000"), -- 41.6 + 76.4 = 118
	(b"11000001110000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100111000000000000000000", b"11000010001011110011001100110011"), -- -24.3 + -19.5 = -43.8
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000010110011001100110", b"11000010101111000110011001100110"), -- 2.5 + -96.7 = -94.2
	(b"11000001100101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111100000000000000000000", b"11000001110100110011001100110011"), -- -18.9 + -7.5 = -26.4
	(b"01000010100100101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011101100000000000000000", b"01000011000001101100110011001101"), -- 73.3 + 61.5 = 134.8
	(b"01000010000100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111001001100110011001101", b"01000010100000110000000000000000"), -- 36.9 + 28.6 = 65.5
	(b"11000010010101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100111001100110011001101", b"11000011000000111110011001100110"), -- -53.5 + -78.4 = -131.9
	(b"01000001101001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001011111001100110011010", b"01000010100000011001100110011010"), -- 20.9 + 43.9 = 64.8
	(b"01000010100101010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000010100000000000000000", b"01000010001000000110011001100110"), -- 74.6 + -34.5 = 40.1
	(b"01000010110001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000010000110011001100110", b"01000010100000001001100110011010"), -- 98.4 + -34.1 = 64.3
	(b"01000010001001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000111001100110011010", b"01000010111101110110011001100111"), -- 41.9 + 81.8 = 123.7
	(b"11000010001101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001011101100110011001101", b"10111111101001100110011001100000"), -- -45 + 43.7 = -1.3
	(b"01000010000100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101001011001100110011010", b"01000010011000111001100110011010"), -- 36.2 + 20.7 = 56.9
	(b"11000010010111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101001000000000000000000", b"11000011000010010001100110011010"), -- -55.1 + -82 = -137.1
	(b"11000010100110110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001010010011001100110011010", b"11000010101101001001100110011001"), -- -77.7 + -12.6 = -90.3
	(b"11000001101010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010011100110011001100110", b"11000010100100100000000000000000"), -- -21.4 + -51.6 = -73
	(b"01000010101001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000011001100110011001101", b"01000010111011000110011001100110"), -- 83 + 35.2 = 118.2
	(b"01000001100001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110000110011001100110", b"11000010100101110000000000000000"), -- 16.7 + -92.2 = -75.5
	(b"11000001111011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001010001100110011001101", b"11000010100100000000000000000000"), -- -29.8 + -42.2 = -72
	(b"01000010101101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101010000000000000000", b"00111110100110011001101000000000"), -- 90.8 + -90.5 = 0.300003
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001001100000000000000000000", b"11000001011011100110011001100110"), -- -3.9 + -11 = -14.9
	(b"01000010101110110000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111111000000000000000000", b"01000010011110000000000000000000"), -- 93.5 + -31.5 = 62
	(b"11000001010111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101000010011001100110011", b"11000010101111010000000000000000"), -- -13.9 + -80.6 = -94.5
	(b"01000010101000110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100110001100110011001101", b"01000000101000110011001100110000"), -- 81.5 + -76.4 = 5.1
	(b"01000001110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001111101011001100110011010", b"11000000110010011001100110011100"), -- 24.4 + -30.7 = -6.3
	(b"01000010000001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111100110011001100110", b"11000010011101110011001100110010"), -- 33.4 + -95.2 = -61.8
	(b"11000001110000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100011110000000000000000", b"01000010001111011001100110011010"), -- -24.1 + 71.5 = 47.4
	(b"11000001110001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100000011100110011001101", b"11000010101100101100110011001101"), -- -24.5 + -64.9 = -89.4
	(b"11000001001110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010110001000011001100110011", b"11000010110110111001100110011001"), -- -11.7 + -98.1 = -109.8
	(b"11000010001110000110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"11000010001000001100110011001100"), -- -46.1 + 5.9 = -40.2
	(b"01000010110001010110011001100110", b"00000000000000000000000000000000"),
	(b"01000001111011100110011001100110", b"01000011000000001000000000000000"), -- 98.7 + 29.8 = 128.5
	(b"11000010100110011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011110100110011001100110", b"11000001011001001100110011010000"), -- -76.9 + 62.6 = -14.3
	(b"11000010001110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001100001011001100110011010", b"11000010011111000000000000000000"), -- -46.3 + -16.7 = -63
	(b"01000010101110010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010110000011001100110011010", b"01000011001111010110011001100110"), -- 92.6 + 96.8 = 189.4
	(b"11000001011001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010111100110011001100110", b"01000010001001010011001100110011"), -- -14.3 + 55.6 = 41.3
	(b"01000010011111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001011001100110011010", b"11000010000011101100110011001110"), -- 63.1 + -98.8 = -35.7
	(b"01000001001010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111100100110011001100110", b"01000010001000111001100110011010"), -- 10.6 + 30.3 = 40.9
	(b"01000010101101001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101011000110011001100110", b"01000000100000110011001101000000"), -- 90.3 + -86.2 = 4.10001
	(b"11000010101001010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110111100110011001100110", b"11000010010110101100110011001101"), -- -82.5 + 27.8 = -54.7
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010001010011001100110011", b"11000010010000111001100110011001"), -- 0.4 + -49.3 = -48.9
	(b"01000010100101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100010010000000000000000", b"01000000111000110011001100110000"), -- 75.6 + -68.5 = 7.1
	(b"01000001010100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001111000000000000000000", b"11000010000001111001100110011010"), -- 13.1 + -47 = -33.9
	(b"01000001101100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100000010110011001100110", b"01000010101011011001100110011001"), -- 22.1 + 64.7 = 86.8
	(b"11000010100011011100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110001011001100110011010", b"11000010001110001100110011001101"), -- -70.9 + 24.7 = -46.2
	(b"01000001101110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001010101001100110011001101", b"01000001000110110011001100110011"), -- 23 + -13.3 = 9.7
	(b"11000010101110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100010100000000000000000", b"11000001101110000000000000000000"), -- -92 + 69 = -23
	(b"11000001001111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000010110011001100110", b"01000010101010011100110011001100"), -- -11.8 + 96.7 = 84.9
	(b"01000001001000110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000001001010110011001100110011"), -- 10.2 + 0.5 = 10.7
	(b"11000010000111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000101101100110011001101", b"11000000000001100110011001100000"), -- -39.8 + 37.7 = -2.1
	(b"11000010101011110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101000000000000000000000", b"11000011001001111000000000000000"), -- -87.5 + -80 = -167.5
	(b"11000010000100010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001110111001100110011010", b"01000001001010011001100110011100"), -- -36.3 + 46.9 = 10.6
	(b"01000001100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010100011001100110011010", b"11000010000100011001100110011010"), -- 16 + -52.4 = -36.4
	(b"11000010100011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110011100110011001100110", b"11000010110000100000000000000000"), -- -71.2 + -25.8 = -97
	(b"01000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010000100000000000000000", b"11000010001110000110011001100110"), -- 2.4 + -48.5 = -46.1
	(b"11000010010111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001010011001100110011", b"11000011000110100011001100110011"), -- -55.6 + -98.6 = -154.2
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000000001110011001100110011010"), -- 0.9 + -3.8 = -2.9
	(b"11000010100000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010001000110011001100110", b"11000010111000110110011001100110"), -- -64.6 + -49.1 = -113.7
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001011101100110011001100110", b"01000001110001100110011001100110"), -- 9.4 + 15.4 = 24.8
	(b"11000010101011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011000010011001100110011", b"11000001111101000000000000000010"), -- -86.8 + 56.3 = -30.5
	(b"11000001110111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011101010011001100110011", b"01000010000001100000000000000000"), -- -27.8 + 61.3 = 33.5
	(b"01000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100110011100110011001101", b"01000001100000001100110011001100"), -- 93 + -76.9 = 16.1
	(b"11000001100010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011001100110011001100110", b"11000010100101010110011001100110"), -- -17.1 + -57.6 = -74.7
	(b"01000010101110101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000010000110011001100110", b"01000010111111101100110011001101"), -- 93.3 + 34.1 = 127.4
	(b"01000000001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000100110011001100110011", b"01000010000111010011001100110011"), -- 2.5 + 36.8 = 39.3
	(b"01000010001011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100001111001100110011010", b"11000001101111110011001100110100"), -- 43.9 + -67.8 = -23.9
	(b"01000010100100010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101000100011001100110011", b"01000011000110011100110011001100"), -- 72.7 + 81.1 = 153.8
	(b"11000010000000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101000000000000000000000", b"11000010010100111001100110011010"), -- -32.9 + -20 = -52.9
	(b"01000001110101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001011001100110011010", b"01000010101110101100110011001101"), -- 26.6 + 66.8 = 93.4
	(b"01000010010110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110101001100110011010", b"11000001101110001100110011001110"), -- 54.2 + -77.3 = -23.1
	(b"01000010100010110011001100110011", b"00000000000000000000000000000000"),
	(b"10000000000000000000000000000000", b"01000010100010110011001100110011"), -- 69.6 + -0 = 69.6
	(b"11000001100101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000001101101011001100110011001"), -- -18.9 + -3.8 = -22.7
	(b"01000001100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101111000000000000000000", b"11000000110010011001100110011000"), -- 17.2 + -23.5 = -6.3
	(b"01000010010111000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000010011111001100110011001100"), -- 55.1 + 8.1 = 63.2
	(b"01000010011101000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000111000000000000000000", b"01000010110010000011001100110011"), -- 61.1 + 39 = 100.1
	(b"11000010010011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100010100110011001100110", b"11000010100010011100110011001100"), -- -51.6 + -17.3 = -68.9
	(b"01000010101011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010001000110011001100110", b"01000011000010001011001100110011"), -- 87.6 + 49.1 = 136.7
	(b"01000001011110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100000011001100110011010", b"11000010010001000110011001100111"), -- 15.7 + -64.8 = -49.1
	(b"11000001101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000110101100110011001101", b"11000010011100101100110011001101"), -- -22 + -38.7 = -60.7
	(b"01000010001001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000110110011001100110", b"01000011000010101100110011001100"), -- 41.1 + 97.7 = 138.8
	(b"11000010000101111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001101001100110011001101", b"01000000111010011001100110011000"), -- -37.9 + 45.2 = 7.3
	(b"01000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100001100110011001100110", b"01000001110101001100110011001100"), -- 9.8 + 16.8 = 26.6
	(b"01000010000100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100110100110011001100110", b"01000001100010100110011001100110"), -- 36.6 + -19.3 = 17.3
	(b"11000001110010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000111000000000000000000", b"01000001011000000000000000000000"), -- -25 + 39 = 14
	(b"11000010101000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001010010110011001100110011", b"11000010100010100011001100110100"), -- -81.8 + 12.7 = -69.1
	(b"11000010000010100000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000010000110001100110011001101"), -- -34.5 + -3.7 = -38.2
	(b"11000010011111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000011100110011001101", b"01000010000001101100110011001101"), -- -63.2 + 96.9 = 33.7
	(b"01000010001001111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100101110000000000000000", b"11000010000001100110011001100110"), -- 41.9 + -75.5 = -33.6
	(b"11000010000001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001100011001100110011010", b"01000001001010110011001100110100"), -- -33.7 + 44.4 = 10.7
	(b"01000010011101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000100100110011001100110", b"01000001110001001100110011001110"), -- 61.2 + -36.6 = 24.6
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101010010000000000000000", b"11000010101010000000000000000000"), -- 0.5 + -84.5 = -84
	(b"01000010101011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111010000000000000000000", b"01000010111010010011001100110011"), -- 87.6 + 29 = 116.6
	(b"11000010100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100011001001100110011010", b"11000011000100100100110011001101"), -- -76 + -70.3 = -146.3
	(b"11000010011110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011011111001100110011010", b"11000000001100110011001100110000"), -- -62.7 + 59.9 = -2.8
	(b"11000010100011000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011100111001100110011010", b"11000001000100110011001100110000"), -- -70.1 + 60.9 = -9.2
	(b"01000010001101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101001001100110011010", b"01000010111100000011001100110100"), -- 45.8 + 74.3 = 120.1
	(b"01000010101000110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100000100000000000000000", b"01000001100001011001100110011000"), -- 81.7 + -65 = 16.7
	(b"01000001010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001011100000000000000000000", b"01000001110110000000000000000000"), -- 12 + 15 = 27
	(b"11000010011111010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001001100110011001100110011", b"11000010100101010000000000000000"), -- -63.3 + -11.2 = -74.5
	(b"11000010101100111100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101110001100110011001101", b"11000010100001011001100110011010"), -- -89.9 + 23.1 = -66.8
	(b"01000010010100010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100111001100110011001101", b"01000011000000101011001100110011"), -- 52.3 + 78.4 = 130.7
	(b"11000010010001011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"11000010001110100110011001100111"), -- -49.4 + 2.8 = -46.6
	(b"01000010000100100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111011011001100110011010", b"01000000110110011001100110011000"), -- 36.5 + -29.7 = 6.8
	(b"01000010101111001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001111001100110011010", b"01000011001100100001100110011010"), -- 94.3 + 83.8 = 178.1
	(b"01000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011010011001100110011010", b"01000010100000000110011001100111"), -- 5.8 + 58.4 = 64.2
	(b"01000010101110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001001010011001100110011010", b"01000010101000111001100110011010"), -- 92.4 + -10.6 = 81.8
	(b"01000010100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001101010000000000000000000", b"01000010110000111001100110011010"), -- 76.8 + 21 = 97.8
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000000110000110011001100110011"), -- -6.2 + 0.1 = -6.1
	(b"11000010101010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001100000000000000000000000", b"11000010100010010011001100110011"), -- -84.6 + 16 = -68.6
	(b"01000010011011101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100000111100110011001101", b"11000000110001100110011001101000"), -- 59.7 + -65.9 = -6.2
	(b"01000010001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100011111100110011001101", b"01000010111000110000000000000000"), -- 41.6 + 71.9 = 113.5
	(b"01000010100010000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101101110000000000000000", b"01000011000111111001100110011010"), -- 68.1 + 91.5 = 159.6
	(b"01000001100110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101110100011001100110011", b"01000010111000001100110011001100"), -- 19.3 + 93.1 = 112.4
	(b"11000010101010110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000100000000000000000000", b"11000010111100110000000000000000"), -- -85.5 + -36 = -121.5
	(b"01000001100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011010011001100110011010", b"01000010100110001100110011001101"), -- 18 + 58.4 = 76.4
	(b"11000010100011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001011010011001100110011", b"11000010111001001001100110011010"), -- -71 + -43.3 = -114.3
	(b"01000010100111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100001010011001100110011", b"01000011000100001001100110011010"), -- 78 + 66.6 = 144.6
	(b"01000001101010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100010000110011001100110", b"01000010101100110000000000000000"), -- 21.3 + 68.2 = 89.5
	(b"01000001101100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100111010110011001100110", b"11000010011000011111111111111111"), -- 22.2 + -78.7 = -56.5
	(b"11000010110000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000011100110011001101", b"11000011001100101011001100110100"), -- -97.8 + -80.9 = -178.7
	(b"01000010100000110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001011010000000000000000000", b"01000010101000000110011001100110"), -- 65.7 + 14.5 = 80.2
	(b"01000010010001011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100111010011001100110011", b"01000011000000000000000000000000"), -- 49.4 + 78.6 = 128
	(b"01000010101011010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000101001100110011001101", b"01000010111101111001100110011010"), -- 86.6 + 37.2 = 123.8
	(b"11000010100110010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000000110011001100110011", b"11000010001011111001100110011001"), -- -76.7 + 32.8 = -43.9
	(b"01000001110111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111101100110011001100110", b"11000000010000000000000000000000"), -- 27.8 + -30.8 = -3
	(b"01000010001110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010001001100110011001101", b"01000010101111101100110011001101"), -- 46.2 + 49.2 = 95.4
	(b"01000010100010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110001110011001100110011", b"01000010101110011100110011001101"), -- 68 + 24.9 = 92.9
	(b"11000010011100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011110111001100110011010", b"01000000000110011001100110100000"), -- -60.5 + 62.9 = 2.4
	(b"01000001110001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001001001100110011001101", b"01000010100001000011001100110011"), -- 24.9 + 41.2 = 66.1
	(b"01000010100111010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100110100000000000000000", b"01000011000110111000000000000000"), -- 78.5 + 77 = 155.5
	(b"01000010001110100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111010011001100110011001101", b"01000010001101110011001100110011"), -- 46.6 + -0.8 = 45.8
	(b"01000010010101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111100110011001100110011", b"01000001101110011001100110011001"), -- 53.6 + -30.4 = 23.2
	(b"01000010010000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"01000010000111001100110011001100"), -- 48.1 + -8.9 = 39.2
	(b"01000010110000110110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"01000010110010110110011001100110"), -- 97.7 + 4 = 101.7
	(b"11000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001100101100110011001101", b"11000010010101001100110011001101"), -- -8.5 + -44.7 = -53.2
	(b"11000001101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001100100000000000000000", b"01000001101101110011001100110011"), -- -21.6 + 44.5 = 22.9
	(b"11000001011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101111100011001100110011", b"01000010100111111100110011001101"), -- -15.2 + 95.1 = 79.9
	(b"01000001110010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010101110011001100110011", b"11000001111001100110011001100110"), -- 25 + -53.8 = -28.8
	(b"11000010100101011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100101101001100110011010", b"00111110110011001100110100000000"), -- -74.9 + 75.3 = 0.400002
	(b"11000001100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101001011001100110011010", b"11000010000111100000000000000000"), -- -18.8 + -20.7 = -39.5
	(b"11000010101100110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011110110011001100110", b"11000011001100010110011001100110"), -- -89.7 + -87.7 = -177.4
	(b"11000010100010111100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111101000000000000000000", b"11000010110010001100110011001101"), -- -69.9 + -30.5 = -100.4
	(b"11000001001100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100001001001100110011010", b"01000010010111010011001100110100"), -- -11 + 66.3 = 55.3
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"10111111111100110011001100110100"), -- 3.5 + -5.4 = -1.9
	(b"11000001111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110010110011001100110", b"11000010110101001001100110011001"), -- -29.6 + -76.7 = -106.3
	(b"01000010000110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111001001100110011001101", b"01000001000110011001100110011010"), -- 38.2 + -28.6 = 9.6
	(b"01000010000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101010110011001100110", b"11000010011000101100110011001100"), -- 34 + -90.7 = -56.7
	(b"11000010110000101001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110101100110011001100110", b"11000010101101010011001100110100"), -- -97.3 + 6.7 = -90.6
	(b"01000010110000011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111000100110011001100110", b"01000010100010010011001100110100"), -- 96.9 + -28.3 = 68.6
	(b"11000010101000010011001100110011", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000010100111101001100110011001"), -- -80.6 + 1.3 = -79.3
	(b"11000001100000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111101001100110011001101", b"11000010001110101100110011001101"), -- -16.1 + -30.6 = -46.7
	(b"01000001101111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011011100110011001100110", b"11000010000100000110011001100110"), -- 23.5 + -59.6 = -36.1
	(b"11000010000101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000100100110011001100110", b"10111111100110011001100110100000"), -- -37.8 + 36.6 = -1.2
	(b"11000010100110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110000011001100110011010", b"11000011001011010000000000000000"), -- -76.2 + -96.8 = -173
	(b"11000010100111011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010000000000000000000000", b"11000010111111011100110011001101"), -- -78.9 + -48 = -126.9
	(b"01000010100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001001000110011001100110", b"01000010111000100011001100110011"), -- 72 + 41.1 = 113.1
	(b"11000010101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101001010000000000000000", b"11000000111000110011001100110000"), -- -89.6 + 82.5 = -7.1
	(b"11000010100101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010110110011001100110", b"11000011000100011000000000000000"), -- -75.8 + -69.7 = -145.5
	(b"01000000110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001101000110011001100110", b"11000010000110010011001100110011"), -- 6.8 + -45.1 = -38.3
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101101000011001100110011", b"01000010110000000110011001100110"), -- 6.1 + 90.1 = 96.2
	(b"01000010100101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001001110011001100110011010", b"01000010011110110011001100110100"), -- 74.4 + -11.6 = 62.8
	(b"01000010101111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011010100110011001100110", b"01000011000110100110011001100110"), -- 95.8 + 58.6 = 154.4
	(b"11000010100110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001001100110011001101", b"11000011001011101001100110011010"), -- -76.2 + -98.4 = -174.6
	(b"11000001010011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001010011001100110011001101", b"10111101110011001100110010000000"), -- -12.9 + 12.8 = -0.0999994
	(b"01000010001010000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100011001100110011001101", b"01000001110000111111111111111111"), -- 42.1 + -17.6 = 24.5
	(b"01000010010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101101011100110011001101", b"11000010000111101100110011001101"), -- 51.2 + -90.9 = -39.7
	(b"01000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100011111100110011001101", b"11000010100010010110011001100111"), -- 3.2 + -71.9 = -68.7
	(b"01000010010111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101101001100110011010", b"11000010000100001100110011001110"), -- 55.1 + -91.3 = -36.2
	(b"11000010011111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101101001001100110011010", b"01000001110101110011001100110100"), -- -63.4 + 90.3 = 26.9
	(b"01000001100110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111000100110011001100110", b"01000010001111101100110011001100"), -- 19.4 + 28.3 = 47.7
	(b"01000010000011101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110011100110011001100110", b"01000001000111100110011001101000"), -- 35.7 + -25.8 = 9.9
	(b"11000010010000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010110011001100110011", b"01000010000100101100110011001100"), -- -48.9 + 85.6 = 36.7
	(b"11000001011010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101011100011001100110011", b"01000010100100001100110011001101"), -- -14.7 + 87.1 = 72.4
	(b"01000010101000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001110000000000000000", b"01000011000100111110011001100110"), -- 80.4 + 67.5 = 147.9
	(b"11000001011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001001011100110011001100110", b"11000001110010100110011001100110"), -- -14.4 + -10.9 = -25.3
	(b"01000010011011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"01000010011110000000000000000000"), -- 59.7 + 2.3 = 62
	(b"01000010101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100111111100110011001101", b"01000011000111111110011001100110"), -- 80 + 79.9 = 159.9
	(b"01000010000110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011001100110011001100110", b"11000001100101011001100110011000"), -- 38.9 + -57.6 = -18.7
	(b"01000010011001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011110011001100110011010", b"01000010111100001001100110011010"), -- 57.9 + 62.4 = 120.3
	(b"11000001101110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000110110011001100110011", b"01000001011110110011001100110010"), -- -23.1 + 38.8 = 15.7
	(b"01000001100110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100111010011001100110011", b"01000010110000110011001100110011"), -- 19 + 78.6 = 97.6
	(b"01000001101100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"01000001100101001100110011001100"), -- 22.3 + -3.7 = 18.6
	(b"11000010100100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000000001110011001100110011010", b"11000010100101100011001100110011"), -- -72.2 + -2.9 = -75.1
	(b"11000010101110010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100100011001100110011010", b"11000001100111100110011001100100"), -- -92.6 + 72.8 = -19.8
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100011101001100110011010", b"11000010100011010000000000000000"), -- 0.8 + -71.3 = -70.5
	(b"01000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000110010011001100110011", b"11000001111100001100110011001100"), -- 8.2 + -38.3 = -30.1
	(b"11000010100100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001001101001100110011001101", b"11000010101010010000000000000000"), -- -73.2 + -11.3 = -84.5
	(b"11000001111010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001000000000000000000000", b"01000001001010011001100110011010"), -- -29.4 + 40 = 10.6
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110010011001100110011001101", b"11000001000010110011001100110011"), -- -8.9 + 0.2 = -8.7
	(b"11000010101101010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011001111001100110011010", b"11000011000101000110011001100110"), -- -90.5 + -57.9 = -148.4
	(b"11000010110001010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101111000000000000000000", b"11000000100101100110011001100000"), -- -98.7 + 94 = -4.7
	(b"11000001001101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110011001100110011001101", b"01000001011000110011001100110100"), -- -11.4 + 25.6 = 14.2
	(b"01000010001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110001010011001100110011", b"01000011000011110000000000000000"), -- 44.4 + 98.6 = 143
	(b"01000010101011001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011010110011001100110011", b"01000011000100010001100110011010"), -- 86.3 + 58.8 = 145.1
	(b"01000010101001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000011000110011001100110", b"01000010111011010110011001100110"), -- 83.6 + 35.1 = 118.7
	(b"11000010011111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011100010011001100110011", b"11000010111110000011001100110011"), -- -63.8 + -60.3 = -124.1
	(b"10111111100011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001111111001100110011010", b"01000010001110110011001100110100"), -- -1.1 + 47.9 = 46.8
	(b"01000001010101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111110011001100110011010", b"01000001101010011001100110011010"), -- 13.4 + 7.8 = 21.2
	(b"01000010010100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001001100110011001100110011", b"01000010011111011001100110011010"), -- 52.2 + 11.2 = 63.4
	(b"01000001001111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100111111001100110011010", b"01000010101101110110011001100111"), -- 11.9 + 79.8 = 91.7
	(b"11000010100100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100101100110011001100110", b"11000010100111010000000000000000"), -- -73.8 + -4.7 = -78.5
	(b"01000010101000010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111011000000000000000000", b"01000010010011000000000000000000"), -- 80.5 + -29.5 = 51
	(b"01000001111100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001110111110011001100110011", b"01000010011010000110011001100110"), -- 30.2 + 27.9 = 58.1
	(b"01000010000010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001100110001100110011001101", b"01000001011100011001100110011010"), -- 34.2 + -19.1 = 15.1
	(b"11000010001101010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000011000110011001100110", b"11000001001000110011001100110100"), -- -45.3 + 35.1 = -10.2
	(b"11000010100110100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010110000000000000000", b"11000000111100110011001100110000"), -- -77.1 + 69.5 = -7.6
	(b"01000001110011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001011010110011001100110011", b"01000010001000011001100110011010"), -- 25.7 + 14.7 = 40.4
	(b"01000010100011010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011001011001100110011010", b"01000001010100011001100110011000"), -- 70.5 + -57.4 = 13.1
	(b"11000010011010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100011100110011001100110", b"11000010100101111001100110011010"), -- -58 + -17.8 = -75.8
	(b"11000010100001000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010110000010011001100110011", b"11000011001000101011001100110011"), -- -66.1 + -96.6 = -162.7
	(b"01000001110100100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000001110100000000000000000000"), -- 26.3 + -0.3 = 26
	(b"11000010101101011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010110111001100110011010", b"11000010000100000000000000000000"), -- -90.9 + 54.9 = -36
	(b"11000010100111111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110001011001100110011010", b"01000001100101110011001100110100"), -- -79.9 + 98.8 = 18.9
	(b"11000010110001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100100100011001100110011", b"11000001110101000000000000000000"), -- -99.6 + 73.1 = -26.5
	(b"11000001101110001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000001101011110011001100110011"), -- -23.1 + 1.2 = -21.9
	(b"01000010101000000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100111000110011001100110", b"00111111111100110011001101000000"), -- 80.1 + -78.2 = 1.9
	(b"11000010101001111001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100011001100110011001101", b"11000010101100000110011001100111"), -- -83.8 + -4.4 = -88.2
	(b"11000010101011110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011111011001100110011010", b"11000011000101110001100110011010"), -- -87.7 + -63.4 = -151.1
	(b"11000010100101111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001111010011001100110011", b"11000010111101100110011001100110"), -- -75.9 + -47.3 = -123.2
	(b"01000010011111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101001001100110011001101", b"01000010101010000011001100110011"), -- 63.5 + 20.6 = 84.1
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001010101100110011001101", b"01000010000010011001100110011010"), -- -8.3 + 42.7 = 34.4
	(b"11000010101100110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001111111001100110011001101", b"11000010011010000110011001100110"), -- -89.7 + 31.6 = -58.1
	(b"11000010110000000011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000010110011001100110011", b"11000010101011101100110011001101"), -- -96.1 + 8.7 = -87.4
	(b"11000010101001100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101001100110011001100110", b"11000011001001100100110011001100"), -- -83.1 + -83.2 = -166.3
	(b"11000010001100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010110001101100110011001101", b"11000011000011111001100110011010"), -- -44.2 + -99.4 = -143.6
	(b"11000010000101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000101000110011001100110", b"10111110110011001100110100000000"), -- -37.5 + 37.1 = -0.400002
	(b"11000010101011100011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111110011001100110011010", b"11000010010111111001100110011001"), -- -87.1 + 31.2 = -55.9
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010011100000000000000000", b"11000010011100110011001100110011"), -- -9.3 + -51.5 = -60.8
	(b"11000010001100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010100110011001100110", b"11000010111001000011001100110011"), -- -44.9 + -69.2 = -114.1
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110111001100110011010", b"11000010101001111100110011001101"), -- -6.1 + -77.8 = -83.9
	(b"01000010001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011100111001100110011010", b"01000010110101101001100110011010"), -- 46.4 + 60.9 = 107.3
	(b"11000001110111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110011100110011001101", b"11000010110100011001100110011010"), -- -27.9 + -76.9 = -104.8
	(b"11000000010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101111000000000000000000", b"01000001101000011001100110011010"), -- -3.3 + 23.5 = 20.2
	(b"01000010011001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010010110011001100110", b"01000010111111010000000000000000"), -- 57.8 + 68.7 = 126.5
	(b"11000010001001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010111111001100110011010", b"11000010110000011100110011001101"), -- -41 + -55.9 = -96.9
	(b"01000010000100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001101111001100110011001101", b"01000001010010011001100110011010"), -- 36.2 + -23.6 = 12.6
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000100000000000000000000", b"01000010001011011001100110011010"), -- 7.4 + 36 = 43.4
	(b"01000010101010010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110010110011001100110011", b"01000010110110111100110011001101"), -- 84.5 + 25.4 = 109.9
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010110001011100110011001101", b"11000010101101110000000000000000"), -- 7.4 + -98.9 = -91.5
	(b"11000010001101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001100011001100110011010", b"10111111000110011001100110000000"), -- -45 + 44.4 = -0.599998
	(b"01000010010101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101011001100110011001101", b"01000011000011000011001100110011"), -- 53.8 + 86.4 = 140.2
	(b"11000010010001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101100100011001100110011", b"01000010001000000000000000000000"), -- -49.1 + 89.1 = 40
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010111100000000000000000", b"11000010010000110011001100110011"), -- 6.7 + -55.5 = -48.8
	(b"11000001101000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111010100110011001100110", b"11000010010001100000000000000000"), -- -20.2 + -29.3 = -49.5
	(b"01000010011111100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000100000000000000000000", b"01000001110111000000000000000000"), -- 63.5 + -36 = 27.5
	(b"11000010100010010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010110100110011001100110", b"11000010111101100110011001100110"), -- -68.6 + -54.6 = -123.2
	(b"11000010011011000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000000111001100110011010", b"11000010101110000000000000000000"), -- -59.1 + -32.9 = -92
	(b"01000010100001011100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110010000000000000000000", b"01000010101101111100110011001101"), -- 66.9 + 25 = 91.9
	(b"01000010000010100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111101100110011001101", b"01000010101101000110011001100110"), -- 34.5 + 55.7 = 90.2
	(b"01000010001010101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101001010011001100110011", b"11000010000111111001100110011001"), -- 42.7 + -82.6 = -39.9
	(b"01000010000010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110100011001100110011010", b"01000001000001100110011001100100"), -- 34.6 + -26.2 = 8.4
	(b"11000001110101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101001010110011001100110", b"11000010110110101100110011001100"), -- -26.7 + -82.7 = -109.4
	(b"11000010000101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010101010011001100110011", b"01000001100000100110011001100110"), -- -37 + 53.3 = 16.3
	(b"01000001010010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000101001100110011001101", b"01000010010001101100110011001101"), -- 12.5 + 37.2 = 49.7
	(b"11000010100011111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100001001001100110011010", b"11000011000010100011001100110100"), -- -71.9 + -66.3 = -138.2
	(b"11000010100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001000000110011001100110", b"11000010111000110110011001100110"), -- -73.6 + -40.1 = -113.7
	(b"11000010100001100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010000100110011001100110", b"11000001100101000000000000000000"), -- -67.1 + 48.6 = -18.5
	(b"11000010100010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011010101100110011001101", b"11000001000101001100110011001100"), -- -68 + 58.7 = -9.3
	(b"01000010100101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000010000000000000000000", b"01000010110110000000000000000000"), -- 74 + 34 = 108
	(b"11000010001110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010000011001100110011", b"01000001101010100110011001100110"), -- -46.8 + 68.1 = 21.3
	(b"11000010101100010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000001001100110011001101", b"11000010111100110110011001100110"), -- -88.5 + -33.2 = -121.7
	(b"01000010101100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101110100110011001100110", b"01000010110111110110011001100110"), -- 88.4 + 23.3 = 111.7
	(b"01000010011111101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001011010011001100110011010", b"01000010100111001001100110011010"), -- 63.7 + 14.6 = 78.3
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101110001001100110011010", b"01000010101001100011001100110100"), -- -9.2 + 92.3 = 83.1
	(b"11000001111111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010111000110011001100110", b"11000010101011010110011001100110"), -- -31.6 + -55.1 = -86.7
	(b"01000010001110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101001100011001100110011", b"01000011000000011001100110011010"), -- 46.5 + 83.1 = 129.6
	(b"01000010001110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100101011100110011001101", b"01000010111100110000000000000000"), -- 46.6 + 74.9 = 121.5
	(b"01000010110001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010100011001100110011010", b"01000011000101111100110011001101"), -- 99.4 + 52.4 = 151.8
	(b"11000010100100011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100000011100110011001101", b"11000001000000000000000000000000"), -- -72.9 + 64.9 = -8
	(b"11000001000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000011100110011001100110", b"11000010001100110011001100110011"), -- -9.2 + -35.6 = -44.8
	(b"11000001110000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011100110011001100110011", b"11000010101010100011001100110011"), -- -24.3 + -60.8 = -85.1
	(b"01000010101100111100110011001101", b"00000000000000000000000000000000"),
	(b"11000001100101000000000000000000", b"01000010100011101100110011001101"), -- 89.9 + -18.5 = 71.4
	(b"11000010010000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011100101100110011001101", b"11000010110110110011001100110100"), -- -48.9 + -60.7 = -109.6
	(b"11000010101110110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010000001100110011001101", b"11000010001101010011001100110011"), -- -93.5 + 48.2 = -45.3
	(b"11000001101010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011110001100110011001101", b"01000010001001001100110011001101"), -- -21 + 62.2 = 41.2
	(b"11000010101010111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101111100000000000000000", b"11000011001101001110011001100110"), -- -85.9 + -95 = -180.9
	(b"11000010100101101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101110010000000000000000", b"01000001100010001100110011001100"), -- -75.4 + 92.5 = 17.1
	(b"01000010101011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100001100000000000000000", b"01000001101001001100110011001100"), -- 87.6 + -67 = 20.6
	(b"01000010100010011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111001110011001100110011", b"01000010001000000000000000000000"), -- 68.9 + -28.9 = 40
	(b"01000010000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010110000000000000000", b"11000010010000101100110011001101"), -- 36.8 + -85.5 = -48.7
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111011001100110011001101", b"11000010000011000000000000000000"), -- -5.4 + -29.6 = -35
	(b"01000010100000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011001001100110011010", b"11000001101011001100110011010000"), -- 64.7 + -86.3 = -21.6
	(b"01000001101111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111110011001100110011", b"11000010100011111100110011001100"), -- 23.7 + -95.6 = -71.9
	(b"01000010011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111000000000000000000", b"01000010110111100000000000000000"), -- 56 + 55 = 111
	(b"11000001100110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001100000110011001100110", b"01000001110001100110011001100110"), -- -19.3 + 44.1 = 24.8
	(b"11000010100101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110101011001100110011010", b"11000010001111101100110011001101"), -- -74.4 + 26.7 = -47.7
	(b"11000010101001101001100110011010", b"00000000000000000000000000000000"),
	(b"11000000000011001100110011001101", b"11000010101010110000000000000000"), -- -83.3 + -2.2 = -85.5
	(b"01000001110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001000000110011001100110", b"01000010100001110110011001100110"), -- 27.6 + 40.1 = 67.7
	(b"01000010100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101010100000000000000000", b"01000011000111010000000000000000"), -- 72 + 85 = 157
	(b"11000000000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110110001100110011001101", b"01000001110001100110011001100111"), -- -2.3 + 27.1 = 24.8
	(b"01000010010101000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001001000110011001100110011", b"01000010001010111001100110011001"), -- 53.1 + -10.2 = 42.9
	(b"11000001011010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010110010011001100110011", b"01000010000111100110011001100110"), -- -14.7 + 54.3 = 39.6
	(b"01000010010101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111100011001100110011010", b"01000001101110100110011001100110"), -- 53.5 + -30.2 = 23.3
	(b"10111111110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100101100000000000000000", b"01000010100100101100110011001101"), -- -1.6 + 75 = 73.4
	(b"11000010011111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001111100110011001101", b"11000011000000101110011001100110"), -- -63 + -67.9 = -130.9
	(b"11000010010011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101100001100110011001101", b"01000010000100100110011001100111"), -- -51.8 + 88.4 = 36.6
	(b"11000010101101000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110001111001100110011010", b"01000001000110011001100110100000"), -- -90.2 + 99.8 = 9.60001
	(b"11000010100110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001100111001100110011010", b"11000001111110001100110011001100"), -- -76 + 44.9 = -31.1
	(b"01000010011111100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110001110110011001100110", b"11000010000100001100110011001100"), -- 63.5 + -99.7 = -36.2
	(b"01000010010010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100111001100110011001101", b"11000001111000000000000000000000"), -- 50.4 + -78.4 = -28
	(b"11000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101011010011001100110011", b"01000010100110100110011001100110"), -- -9.4 + 86.6 = 77.2
	(b"01000001110001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010001100000000000000000", b"11000001110001100110011001100110"), -- 24.7 + -49.5 = -24.8
	(b"01000010100010101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101111000110011001100110", b"11000001110001100110011001100100"), -- 69.4 + -94.2 = -24.8
	(b"01000010110001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101110000000000000000000", b"01000000110100110011001100110000"), -- 98.6 + -92 = 6.6
	(b"11000010000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010110010011001100110011", b"01000001011010110011001100110100"), -- -39.6 + 54.3 = 14.7
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000100100110011001100110", b"01000010000100101100110011001100"), -- 0.1 + 36.6 = 36.7
	(b"11000001110110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101100000000000000000000", b"01000010011100111001100110011010"), -- -27.1 + 88 = 60.9
	(b"11000010001100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101010000000000000000", b"11000011000001110110011001100110"), -- -44.9 + -90.5 = -135.4
	(b"11000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001011000000000000000000000", b"01000001000101100110011001100110"), -- -4.6 + 14 = 9.4
	(b"11000010100111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010011100110011001100110", b"11000001110110110011001100110100"), -- -79 + 51.6 = -27.4
	(b"11000010101001001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011111100110011001100110", b"11000001100101011001100110011100"), -- -82.3 + 63.6 = -18.7
	(b"11000001110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001010000000000000000000000", b"11000001011000000000000000000000"), -- -26 + 12 = -14
	(b"11000001101001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011001001100110011010", b"01000010100000110110011001100111"), -- -20.6 + 86.3 = 65.7
	(b"01000010101100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110000011001100110011010", b"01000010100000010011001100110100"), -- 88.8 + -24.2 = 64.6
	(b"01000010010010101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101000101100110011001101", b"01000011000001000001100110011010"), -- 50.7 + 81.4 = 132.1
	(b"11000000100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110000011001100110011010", b"11000001111001011001100110011010"), -- -4.5 + -24.2 = -28.7
	(b"01000010000011000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101000011100110011001101", b"11000010001101111001100110011010"), -- 35 + -80.9 = -45.9
	(b"01000001111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001111100000000000000000", b"01000010100101111100110011001101"), -- 28.4 + 47.5 = 75.9
	(b"11000010011110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000001100000000000000000", b"11000010101111110110011001100110"), -- -62.2 + -33.5 = -95.7
	(b"01000001010001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011001100110011001101", b"01000010110001010110011001100111"), -- 12.3 + 86.4 = 98.7
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011010000000000000000000", b"11000010100000100000000000000000"), -- -7 + -58 = -65
	(b"11000010000011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010010000000000000000", b"11000010111011111100110011001101"), -- -35.4 + -84.5 = -119.9
	(b"11000010100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000110000110011001100110", b"11000010000101000110011001100110"), -- -75.2 + 38.1 = -37.1
	(b"11000010100000100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111111110011001100110011", b"11000010110000011100110011001101"), -- -65 + -31.9 = -96.9
	(b"11000010100000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111110100110011001100110", b"11000010000010001100110011001101"), -- -65.5 + 31.3 = -34.2
	(b"11000001101011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101111010011001100110011", b"01000010100100100011001100110011"), -- -21.5 + 94.6 = 73.1
	(b"01000010101011110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001011001100110011010", b"01000001101001011001100110011000"), -- 87.5 + -66.8 = 20.7
	(b"01000010010100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110111100110011001100110", b"01000001110010001100110011001110"), -- 52.9 + -27.8 = 25.1
	(b"01000010011000100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011000110011001100110011", b"10111110100110011001100110000000"), -- 56.5 + -56.8 = -0.299999
	(b"11000010100101010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100110101100110011001101", b"01000000001110011001100110100000"), -- -74.5 + 77.4 = 2.9
	(b"01000010100000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101100110110011001100110", b"11000001101111110011001100110000"), -- 65.8 + -89.7 = -23.9
	(b"11000010001001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010111010011001100110011", b"01000001010110011001100110011000"), -- -41.7 + 55.3 = 13.6
	(b"01000010000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000101011001100110011010", b"00111110010011001100110000000000"), -- 37.6 + -37.4 = 0.199997
	(b"01000010100010111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000001001100110011010", b"11000001001001100110011001101000"), -- 69.9 + -80.3 = -10.4
	(b"01000010101111010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101110110011001100110", b"01000011001010100100110011001100"), -- 94.6 + 75.7 = 170.3
	(b"01000001010110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010101000110011001100110", b"11000010000111011001100110011001"), -- 13.7 + -53.1 = -39.4
	(b"11000010110001111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010110011001100110011010", b"11000011000110100100110011001101"), -- -99.9 + -54.4 = -154.3
	(b"01000010000001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110010000000000000000000", b"01000010011010010011001100110011"), -- 33.3 + 25 = 58.3
	(b"11000010001100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001101000000000000000000000", b"11000001110001001100110011001100"), -- -44.6 + 20 = -24.6
	(b"01000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001011101100110011001100110", b"11000000101110011001100110011000"), -- 9.6 + -15.4 = -5.8
	(b"11000010001010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010011101100110011001101", b"11000010101111010000000000000000"), -- -42.8 + -51.7 = -94.5
	(b"01000010101001001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001000000110011001100110", b"01000010001010001100110011001110"), -- 82.3 + -40.1 = 42.2
	(b"11000010010100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101000111001100110011010", b"11000011000001011100110011001101"), -- -52 + -81.8 = -133.8
	(b"11000010001101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100100011001100110011010", b"11000010111011010110011001100111"), -- -45.9 + -72.8 = -118.7
	(b"11000010110000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000101100110011001100110", b"11000011000001100100110011001100"), -- -96.7 + -37.6 = -134.3
	(b"01000010110000001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011010111001100110011010", b"01000010000101011001100110011010"), -- 96.3 + -58.9 = 37.4
	(b"01000001100101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110110110011001100110011", b"11000001000011001100110011001100"), -- 18.6 + -27.4 = -8.8
	(b"11000001100111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000100000000000000000", b"01000010011101010011001100110011"), -- -19.7 + 81 = 61.3
	(b"01000010101011001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100001101001100110011010", b"01000011000110011001100110011010"), -- 86.3 + 67.3 = 153.6
	(b"11000010100011111100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110111001100110011001101", b"11000010001100010011001100110100"), -- -71.9 + 27.6 = -44.3
	(b"11000010000000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110001010011001100110011", b"01000010100000111100110011001100"), -- -32.7 + 98.6 = 65.9
	(b"11000001111011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"11000010000011000110011001100110"), -- -29.8 + -5.3 = -35.1
	(b"01000010101111000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001001101100110011001101", b"01000010010100011001100110011001"), -- 94.1 + -41.7 = 52.4
	(b"11000010000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000011011001100110011001101", b"11000010000111101100110011001101"), -- -36 + -3.7 = -39.7
	(b"01000010011000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101011001100110011001101", b"01000011000011101100110011001101"), -- 56.4 + 86.4 = 142.8
	(b"01000010100011011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000011100000000000000000", b"01000010000011011001100110011010"), -- 70.9 + -35.5 = 35.4
	(b"11000001111010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"11000010000011110011001100110011"), -- -29.3 + -6.5 = -35.8
	(b"01000010110000111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100001000000000000000000", b"01000001111111110011001100110100"), -- 97.9 + -66 = 31.9
	(b"11000010101011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111001001100110011010", b"11000011001101100001100110011010"), -- -87.8 + -94.3 = -182.1
	(b"01000010010101000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101110010110011001100110", b"01000011000100011100110011001100"), -- 53.1 + 92.7 = 145.8
	(b"11000010100100001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001011100000000000000000", b"11000010111001111001100110011010"), -- -72.3 + -43.5 = -115.8
	(b"10000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101110110110011001100110", b"01000010101110110110011001100110"), -- -0 + 93.7 = 93.7
	(b"11000010001110111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110000101100110011001101", b"01000010010010100000000000000000"), -- -46.9 + 97.4 = 50.5
	(b"01000001100100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000111001100110011001101", b"01000001111000001100110011001100"), -- 18.3 + 9.8 = 28.1
	(b"01000001100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100000000110011001100110", b"01000010101001100000000000000000"), -- 18.8 + 64.2 = 83
	(b"11000010101011101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010101111001100110011010", b"11000010000001011001100110011010"), -- -87.3 + 53.9 = -33.4
	(b"11000010001101010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101011001001100110011010", b"01000010001001000000000000000001"), -- -45.3 + 86.3 = 41
	(b"01000010100001110000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110010000000000000000000", b"01000010001010100000000000000000"), -- 67.5 + -25 = 42.5
	(b"11000001100100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110110001100110011001101", b"01000001000011001100110011001110"), -- -18.3 + 27.1 = 8.8
	(b"01000010000110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100000111100110011001101", b"11000001110110100110011001101000"), -- 38.6 + -65.9 = -27.3
	(b"01000010100100100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110100000000000000000", b"11000000011110011001100110100000"), -- 73.1 + -77 = -3.9
	(b"01000010010100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001111000110011001100110", b"01000010110001110011001100110011"), -- 52.5 + 47.1 = 99.6
	(b"11000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000001101100110011001101", b"01000001110101100110011001100111"), -- -6.9 + 33.7 = 26.8
	(b"01000010000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100001111100110011001101", b"01000010110101001001100110011010"), -- 38.4 + 67.9 = 106.3
	(b"01000001111100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001111000001100110011001101", b"01000010011010011001100110011010"), -- 30.3 + 28.1 = 58.4
	(b"11000001110100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001100001100110011001101", b"01000001100011100110011001100111"), -- -26.4 + 44.2 = 17.8
	(b"01000001101010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000001101100110011001101", b"01000010010110101100110011001101"), -- 21 + 33.7 = 54.7
	(b"01000010001001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101000011001100110011010", b"01000001101011001100110011001100"), -- 41.8 + -20.2 = 21.6
	(b"01000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011101110011001100110011", b"11000010010110000000000000000000"), -- 7.8 + -61.8 = -54
	(b"11000010000011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001011010011001100110011", b"01000000111100110011001100110000"), -- -35.7 + 43.3 = 7.6
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001001000000000000000000", b"11000010010010111001100110011010"), -- -9.9 + -41 = -50.9
	(b"01000010101101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001011100000000000000000000", b"01000010110101000000000000000000"), -- 91 + 15 = 106
	(b"01000010000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000110011001100110011010", b"01000010001100000000000000000000"), -- 34.4 + 9.6 = 44
	(b"01000001011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100101001001100110011010", b"01000010101100111100110011001101"), -- 15.6 + 74.3 = 89.9
	(b"11000010110001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"11000010101111011100110011001101"), -- -99.8 + 4.9 = -94.9
	(b"01000010001101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000110111001100110011010", b"01000010101010010000000000000000"), -- 45.6 + 38.9 = 84.5
	(b"01000010101101100011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101001100110011001100110", b"01000010101010111100110011001101"), -- 91.1 + -5.2 = 85.9
	(b"01000001011011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011000101100110011001101", b"01000010100011110011001100110011"), -- 14.9 + 56.7 = 71.6
	(b"01000000111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101100100011001100110011", b"01000010110000001001100110011001"), -- 7.2 + 89.1 = 96.3
	(b"01000010100001010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001100110011001100110011", b"01000001101011110011001100110010"), -- 66.7 + -44.8 = 21.9
	(b"01000010000000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"01000001111011100110011001100111"), -- 32.2 + -2.4 = 29.8
	(b"01000010000101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001010101100110011001101", b"11000000101101100110011001101000"), -- 37 + -42.7 = -5.7
	(b"11000010010110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100001010011001100110011", b"11000010111100100110011001100110"), -- -54.6 + -66.6 = -121.2
	(b"01000010101000100011001100110011", b"00000000000000000000000000000000"),
	(b"11000001001010000000000000000000", b"01000010100011010011001100110011"), -- 81.1 + -10.5 = 70.6
	(b"01000010100011010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001011001100110011001101", b"01000010111000110110011001100110"), -- 70.5 + 43.2 = 113.7
	(b"11000010100000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100000100011001100110011", b"10111111001100110011001110000000"), -- -65.8 + 65.1 = -0.700005
	(b"11000010010001111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000001011001100110011010", b"11000010101001101001100110011010"), -- -49.9 + -33.4 = -83.3
	(b"01000010100010101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000110000000000000000", b"01000011001001101110011001100110"), -- 69.4 + 97.5 = 166.9
	(b"11000010010101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000001001100110011001101", b"11000001101001001100110011001100"), -- -53.8 + 33.2 = -20.6
	(b"11000010011111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000010100011001001100110011001"), -- -63.6 + -6.7 = -70.3
	(b"01000010100000001001100110011010", b"00000000000000000000000000000000"),
	(b"01000001010000000000000000000000", b"01000010100110001001100110011010"), -- 64.3 + 12 = 76.3
	(b"11000010100001011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011010110011001100110011", b"11000001000000011001100110011100"), -- -66.9 + 58.8 = -8.1
	(b"01000010100101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100100100011001100110011", b"00111111110110011001100111000000"), -- 74.8 + -73.1 = 1.7
	(b"01000010101001001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011000100000000000000000", b"01000001110011100110011001101000"), -- 82.3 + -56.5 = 25.8
	(b"11000010101111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001011010011001100110011010", b"11000010101000100110011001100111"), -- -95.8 + 14.6 = -81.2
	(b"11000010100101110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010110111001100110011010", b"11000001101001100110011001100100"), -- -75.7 + 54.9 = -20.8
	(b"11000001111110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011110000000000000000000", b"01000001111101011001100110011010"), -- -31.3 + 62 = 30.7
	(b"11000000010011001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100110011001100110011010", b"11000000100011001100110011001101"), -- -3.2 + -1.2 = -4.4
	(b"01000010101110010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101111000110011001100110", b"10111111110110011001100110000000"), -- 92.5 + -94.2 = -1.7
	(b"01000010101011101001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000010110000000011001100110100"), -- 87.3 + 8.8 = 96.1
	(b"01000010101110011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001110110011001100110", b"01000011001000001001100110011010"), -- 92.9 + 67.7 = 160.6
	(b"01000010010110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010110110011001100110011", b"10111111010011001100110011000000"), -- 54 + -54.8 = -0.799999
	(b"11000010101101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"11000010101010000000000000000000"), -- -91 + 7 = -84
	(b"11000010100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000000000110011001100110", b"11000010000001100000000000000000"), -- -65.6 + 32.1 = -33.5
	(b"11000001110100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101001010011001100110011", b"11000010110110011001100110011010"), -- -26.2 + -82.6 = -108.8
	(b"01000010010101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001101001001100110011001101", b"01000010100101000000000000000000"), -- 53.4 + 20.6 = 74
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001000110011001100110011", b"01000010001110000110011001100110"), -- 5.3 + 40.8 = 46.1
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000000100010011001100110011001"), -- -5.7 + 1.4 = -4.3
	(b"01000010000100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000001001100110011010", b"11000010001011111001100110011010"), -- 36.4 + -80.3 = -43.9
	(b"01000010110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001010100110011001100110", b"01000011000011011100110011001100"), -- 99.2 + 42.6 = 141.8
	(b"11000010001001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100100100110011001100110", b"11000010111001000110011001100110"), -- -41 + -73.2 = -114.2
	(b"11000010100111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001110110011001100110011", b"11000010000000001100110011001101"), -- -79 + 46.8 = -32.2
	(b"11000010100110110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101100000011001100110011", b"01000001001001100110011001101000"), -- -77.7 + 88.1 = 10.4
	(b"01000010101010110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110111110011001100110011", b"01000010111000110011001100110011"), -- 85.7 + 27.9 = 113.6
	(b"01000010101100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000011100110011001100110", b"01000010100111111100110011001101"), -- 88.8 + -8.9 = 79.9
	(b"01000010100000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011000011001100110011", b"11000001101001110011001100110100"), -- 65.2 + -86.1 = -20.9
	(b"01000010101101011100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100111110011001100110011", b"01000010110111011001100110011010"), -- 90.9 + 19.9 = 110.8
	(b"11000010101111011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110110110011001100110011", b"11000010111101001001100110011010"), -- -94.9 + -27.4 = -122.3
	(b"01000010001001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101101011001100110011010", b"11000010010001100000000000000001"), -- 41.3 + -90.8 = -49.5
	(b"11000010001010000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110011100110011001100110", b"11000001100000100110011001100110"), -- -42.1 + 25.8 = -16.3
	(b"01000001001000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110100110011001100110011", b"11000001100000100110011001100110"), -- 10.1 + -26.4 = -16.3
	(b"01000010000000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100000011001100110011010", b"11000010000000100000000000000001"), -- 32.3 + -64.8 = -32.5
	(b"11000010000111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100000010011001100110011", b"01000001110011001100110011001100"), -- -39 + 64.6 = 25.6
	(b"01000010110000110110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000010110010101001100110011001"), -- 97.7 + 3.6 = 101.3
	(b"11000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100001100011001100110011", b"11000010100100011001100110011001"), -- -5.7 + -67.1 = -72.8
	(b"01000010101100100011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001100110011001100110011", b"01000010101011001001100110011001"), -- 89.1 + -2.8 = 86.3
	(b"11000010010010100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010101011001100110011010", b"01000000001110011001100110100000"), -- -50.5 + 53.4 = 2.9
	(b"01000010100110100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001001100110011001100110", b"01000010000011011001100110011010"), -- 77 + -41.6 = 35.4
	(b"01000010100101110000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000010100110110110011001100110"), -- 75.5 + 2.2 = 77.7
	(b"01000010100101011100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"01000010100010001001100110011010"), -- 74.9 + -6.6 = 68.3
	(b"11000010101011100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101111101100110011001101", b"01000001000001001100110011010000"), -- -87.1 + 95.4 = 8.3
	(b"11000010001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101011011100110011001101", b"01000010001010100000000000000000"), -- -44.4 + 86.9 = 42.5
	(b"11000010001010110011001100110011", b"00000000000000000000000000000000"),
	(b"00111111010011001100110011001101", b"11000010001010000000000000000000"), -- -42.8 + 0.8 = -42
	(b"01000001100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000000011001100110011010", b"01000001000010110011001100110010"), -- 16.8 + -8.1 = 8.7
	(b"01000010010100010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100011010011001100110011", b"11000001100100100110011001100110"), -- 52.3 + -70.6 = -18.3
	(b"11000010000111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001001111001100110011010", b"11000010101000110110011001100110"), -- -39.8 + -41.9 = -81.7
	(b"01000010100100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001101100110011001100110", b"01000010111010110011001100110011"), -- 72 + 45.6 = 117.6
	(b"11000010011110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101100010011001100110011", b"11000011000101110110011001100110"), -- -62.8 + -88.6 = -151.4
	(b"01000010001110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011100001100110011001101", b"01000010110101100000000000000000"), -- 46.8 + 60.2 = 107
	(b"01000010101010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100111111100110011001101", b"01000000100100000000000000000000"), -- 84.4 + -79.9 = 4.5
	(b"01000010001101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100011011001100110011010", b"01000010011110111001100110011010"), -- 45.2 + 17.7 = 62.9
	(b"11000010100001011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101111000011001100110011", b"01000001110110011001100110011000"), -- -66.9 + 94.1 = 27.2
	(b"11000010100101110000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100100100110011001100110", b"11000010101110111001100110011010"), -- -75.5 + -18.3 = -93.8
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100001000000000000000000", b"01000000111001100110011001100110"), -- -9.3 + 16.5 = 7.2
	(b"11000001001110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000000100000000000000000", b"11000010001100001100110011001101"), -- -11.7 + -32.5 = -44.2
	(b"01000010010000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"01000010000111000000000000000000"), -- 48.7 + -9.7 = 39
	(b"11000010000010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000010001100101100110011001101"), -- -34.9 + -9.8 = -44.7
	(b"11000010001111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001010001100110011001101", b"11000010101100111001100110011010"), -- -47.6 + -42.2 = -89.8
	(b"11000010000101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001010100011001100110011010", b"11000010010011000000000000000000"), -- -37.9 + -13.1 = -51
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000101011001100110011010", b"01000010001011100000000000000000"), -- 6.1 + 37.4 = 43.5
	(b"01000001111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011101000110011001100110", b"11000010000000010011001100110011"), -- 28.8 + -61.1 = -32.3
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101100011001100110011010", b"01000010101000010000000000000000"), -- -8.3 + 88.8 = 80.5
	(b"11000010100010100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100101110011001100110011", b"11000011000100001001100110011010"), -- -69 + -75.6 = -144.6
	(b"01000010100101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010010111001100110011010", b"01000010111110101001100110011010"), -- 74.4 + 50.9 = 125.3
	(b"11000001100011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100111100110011001100110", b"11000010110000100011001100110011"), -- -17.9 + -79.2 = -97.1
	(b"01000010100111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000010011001100110011", b"01000001101110001100110011001110"), -- 79.4 + -56.3 = 23.1
	(b"11000010011111000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101000010011001100110011", b"01000001100011000000000000000000"), -- -63.1 + 80.6 = 17.5
	(b"01000010101000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010100000110011001100110", b"01000011000001011001100110011010"), -- 81.5 + 52.1 = 133.6
	(b"11000010001101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100111100011001100110011", b"11000010111110010110011001100110"), -- -45.6 + -79.1 = -124.7
	(b"01000001010111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001000111001100110011010", b"11000001110110000000000000000001"), -- 13.9 + -40.9 = -27
	(b"01000010010111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000111000000000000000000", b"01000001100000011001100110011010"), -- 55.2 + -39 = 16.2
	(b"11000001111011110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000001111111011001100110011001"), -- -29.9 + -1.8 = -31.7
	(b"01000001011011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011110110011001100110011", b"10111111010011001100110011010000"), -- 14.9 + -15.7 = -0.8
	(b"01000010100011110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011000110011001100110", b"00111111110000000000000000000000"), -- 71.7 + -70.2 = 1.5
	(b"11000010000110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011010111001100110011010", b"01000001101001011001100110011010"), -- -38.2 + 58.9 = 20.7
	(b"11000010011100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101001100110011001101", b"01000001010110011001100110011100"), -- -60.8 + 74.4 = 13.6
	(b"11000010001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000101010011001100110011", b"11000010100110101001100110011010"), -- -40 + -37.3 = -77.3
	(b"11000010101011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000011110011001100110011", b"11000010111101101100110011001100"), -- -87.6 + -35.8 = -123.4
	(b"01000010101100010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001101011011001100110011010", b"01000010100001011001100110011010"), -- 88.5 + -21.7 = 66.8
	(b"01000010010010101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101001100110011001101", b"01000010101111111100110011001101"), -- 50.7 + 45.2 = 95.9
	(b"11000010100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000001011001100110011010", b"11000010110111111001100110011010"), -- -78.4 + -33.4 = -111.8
	(b"11000010101100100011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000010110000101100110011001101"), -- -89.1 + -8.3 = -97.4
	(b"01000010011011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"01000010010110000110011001100111"), -- 59.9 + -5.8 = 54.1
	(b"11000010101001001001100110011010", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000010101001110011001100110100"), -- -82.3 + -1.3 = -83.6
	(b"11000010000101010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001100001110011001100110011", b"11000010010110001100110011001100"), -- -37.3 + -16.9 = -54.2
	(b"11000001010001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001110000000000000000000", b"11000010011010011001100110011010"), -- -12.4 + -46 = -58.4
	(b"11000001011111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100000111001100110011010", b"11000010101000110011001100110100"), -- -15.8 + -65.8 = -81.6
	(b"11000010010111100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111110000000000000000000000", b"11000010011001000110011001100110"), -- -55.6 + -1.5 = -57.1
	(b"11000001010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011100011001100110011010", b"01000010001110110011001100110100"), -- -13.6 + 60.4 = 46.8
	(b"11000010110000000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000100011001100110011010", b"11000011000001001000000000000000"), -- -96.1 + -36.4 = -132.5
	(b"01000010101101110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001101011011001100110011010", b"01000010111000101100110011001100"), -- 91.7 + 21.7 = 113.4
	(b"01000010100010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011110101100110011001101", b"01000011000000110100110011001101"), -- 68.6 + 62.7 = 131.3
	(b"01000001101100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001001011001100110011010", b"01000010011111100000000000000000"), -- 22.1 + 41.4 = 63.5
	(b"11000010010011111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101100001100110011001101", b"01000010000100100000000000000000"), -- -51.9 + 88.4 = 36.5
	(b"01000010001101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100110000011001100110011", b"01000010111100110000000000000000"), -- 45.4 + 76.1 = 121.5
	(b"11000001110001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001101011100110011001100110", b"11000010001110010011001100110011"), -- -24.5 + -21.8 = -46.3
	(b"01000010101000100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100010111001100110011010", b"01000011000101110000000000000000"), -- 81.2 + 69.8 = 151
	(b"11000010100100110000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100101110011001100110011", b"11000010010110100110011001100110"), -- -73.5 + 18.9 = -54.6
	(b"11000010001001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101011001100110011001101", b"11000010111111110110011001100110"), -- -41.3 + -86.4 = -127.7
	(b"11000001101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010011011001100110011010", b"11000010100100101100110011001101"), -- -22 + -51.4 = -73.4
	(b"11000001001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010101001100110011001101", b"11000010011111100110011001100110"), -- -10.4 + -53.2 = -63.6
	(b"01000010000011100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011111000110011001100110", b"01000010110001010011001100110011"), -- 35.5 + 63.1 = 98.6
	(b"11000010011010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001101100011001100110011010", b"11000010000100001100110011001101"), -- -58.4 + 22.2 = -36.2
	(b"01000001010110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011110000110011001100110", b"01000010100101111001100110011001"), -- 13.7 + 62.1 = 75.8
	(b"01000010101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001111011001100110011010", b"01000010001101011001100110011010"), -- 92.8 + -47.4 = 45.4
	(b"11000010110000011100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110111001100110011001101", b"11000010101101000000000000000000"), -- -96.9 + 6.9 = -90
	(b"01000010001111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000010011001100110011", b"11000001000100011001100110011000"), -- 47.2 + -56.3 = -9.1
	(b"11000010000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101100100000000000000000", b"11000010111101100000000000000000"), -- -34 + -89 = -123
	(b"11000010010111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001010110000000000000000000", b"11000010100010100110011001100110"), -- -55.7 + -13.5 = -69.2
	(b"01000001001100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000010100110011001100110", b"01000010001101100110011001100110"), -- 11 + 34.6 = 45.6
	(b"11000010110000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010010000110011001100110", b"11000011000100101110011001100110"), -- -96.8 + -50.1 = -146.9
	(b"11000001000111001100110011001101", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000001001110011001100110011010"), -- -9.8 + -1.8 = -11.6
	(b"01000010100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100111111100110011001101", b"11000001010010110011001100111000"), -- 67.2 + -79.9 = -12.7
	(b"01000001001011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101110110011001100110", b"01000010110011010011001100110011"), -- 10.9 + 91.7 = 102.6
	(b"01000010001101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010001100110011001101", b"11000010000111000000000000000000"), -- 45.4 + -84.4 = -39
	(b"01000010100000011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101010111100110011001101", b"01000011000101101100110011001101"), -- 64.9 + 85.9 = 150.8
	(b"01000001001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010000111001100110011010", b"01000010011010111001100110011010"), -- 10 + 48.9 = 58.9
	(b"01000010000011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111010011001100110011010", b"01000010100000000110011001100110"), -- 35 + 29.2 = 64.2
	(b"01000010101100000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001010000011001100110011010", b"01000010110010001001100110011001"), -- 88.2 + 12.1 = 100.3
	(b"11000010001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100000001001100110011010", b"01000001100011110011001100110100"), -- -46.4 + 64.3 = 17.9
	(b"11000001101010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000011011001100110011010", b"01000001011000000000000000000010"), -- -21.4 + 35.4 = 14
	(b"11000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111101100110011001101", b"11000010000101010011001100110011"), -- -93 + 55.7 = -37.3
	(b"11000001111000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110100110011001100110011", b"11000010000010110011001100110011"), -- -28.2 + -6.6 = -34.8
	(b"10111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101010011100110011001101", b"01000010101010010000000000000000"), -- -0.4 + 84.9 = 84.5
	(b"01000001101101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100000110011001100110", b"11000010010001010011001100110010"), -- 22.9 + -72.2 = -49.3
	(b"01000010001000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100010100000000000000000", b"01000010110110101100110011001101"), -- 40.4 + 69 = 109.4
	(b"01000010000100100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100101001100110011001101", b"01000001100011110011001100110011"), -- 36.5 + -18.6 = 17.9
	(b"11000010101100010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100111010000000000000000", b"11000011001001110000000000000000"), -- -88.5 + -78.5 = -167
	(b"01000010101110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100011111100110011001101", b"01000011001000111110011001100110"), -- 92 + 71.9 = 163.9
	(b"11000010100100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100001110011001100110011", b"11000010011000111001100110011010"), -- -73.8 + 16.9 = -56.9
	(b"01000010100101100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010111110011001100110011", b"01000011000000101110011001100110"), -- 75.1 + 55.8 = 130.9
	(b"01000010010001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010111001100110011001101", b"01000010110100011100110011001101"), -- 49.7 + 55.2 = 104.9
	(b"01000010100000010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001100110011001100110011", b"01000001100111011001100110011010"), -- 64.5 + -44.8 = 19.7
	(b"01000001111111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000011100110011001101", b"01000011000000001011001100110011"), -- 31.8 + 96.9 = 128.7
	(b"01000010100000010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010010111001100110011010", b"01000010111001101100110011001101"), -- 64.5 + 50.9 = 115.4
	(b"01000010001000010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101010011001100110011", b"01000010111001011100110011001100"), -- 40.3 + 74.6 = 114.9
	(b"11000010100111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001011101100110011001101", b"11000010111100111100110011001100"), -- -78.2 + -43.7 = -121.9
	(b"11000001011010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011110000110011001100110", b"11000010100110011001100110011001"), -- -14.7 + -62.1 = -76.8
	(b"01000010100010000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001010100000000000000000", b"01000010110111010110011001100110"), -- 68.2 + 42.5 = 110.7
	(b"11000010100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011000101100110011001101", b"11000001010000011001100110011100"), -- -68.8 + 56.7 = -12.1
	(b"11000010101011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010001100110011001100110", b"11000010000101100110011001100110"), -- -87.2 + 49.6 = -37.6
	(b"11000010011010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001001010011001100110011", b"11000001100011000000000000000000"), -- -58.8 + 41.3 = -17.5
	(b"11000010101000000011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000010100111110011001100110011"), -- -80.1 + 0.5 = -79.6
	(b"01000010100001010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000111100110011001101", b"11000001111110110011001100110100"), -- 66.5 + -97.9 = -31.4
	(b"11000000101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000001000100011001100110011010"), -- -5.8 + -3.3 = -9.1
	(b"11000001110111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110100000000000000000", b"01000010010001000110011001100110"), -- -27.9 + 77 = 49.1
	(b"01000001101001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011111010011001100110011", b"11000010001010101100110011001100"), -- 20.6 + -63.3 = -42.7
	(b"01000010011100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010001010011001100110011", b"01000001001011100110011001101000"), -- 60.2 + -49.3 = 10.9
	(b"10111111101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000110000110011001100110", b"01000010000100101100110011001100"), -- -1.4 + 38.1 = 36.7
	(b"11000010101110011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000011011001100110011010", b"11000011000000000100110011001101"), -- -92.9 + -35.4 = -128.3
	(b"01000010100101111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100010110000000000000000", b"01000000110011001100110011010000"), -- 75.9 + -69.5 = 6.4
	(b"11000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011110111001100110011010", b"11000010100010110011001100110011"), -- -6.7 + -62.9 = -69.6
	(b"11000010010011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000001100110011001100110011", b"11000010010000110011001100110011"), -- -51.6 + 2.8 = -48.8
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010011000110011001100110", b"11000010001101101100110011001100"), -- 5.4 + -51.1 = -45.7
	(b"01000010100100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000000100000000000000000", b"01000010001000101100110011001100"), -- 73.2 + -32.5 = 40.7
	(b"11000001010000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011110100110011001100110", b"11000010100101010110011001100110"), -- -12.1 + -62.6 = -74.7
	(b"11000001111001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001100011001100110011010", b"11000010100100100011001100110100"), -- -28.7 + -44.4 = -73.1
	(b"01000010100001010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101001001100110011001101", b"01000010001110000110011001100110"), -- 66.7 + -20.6 = 46.1
	(b"01000010000111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110000000000000000000", b"11000010010100100110011001100110"), -- 39.4 + -92 = -52.6
	(b"11000010110001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"11000010101111010011001100110011"), -- -98.2 + 3.6 = -94.6
	(b"11000010100101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000011111001100110011010", b"11000010110111110000000000000000"), -- -75.6 + -35.9 = -111.5
	(b"11000010011001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001001001100110011001100110", b"11000010100001101100110011001101"), -- -57 + -10.4 = -67.4
	(b"01000010110001011100110011001101", b"00000000000000000000000000000000"),
	(b"10111110100110011001100110011010", b"01000010110001010011001100110011"), -- 98.9 + -0.3 = 98.6
	(b"01000010010101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001110101100110011001101", b"01000000110010011001100110011000"), -- 53 + -46.7 = 6.3
	(b"11000001110101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000011001100110011010", b"11000010111101101001100110011010"), -- -26.5 + -96.8 = -123.3
	(b"01000001110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100000110000000000000000", b"11000010001001100000000000000000"), -- 24 + -65.5 = -41.5
	(b"11000010010101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011101100110011001101", b"11000011000011000110011001100110"), -- -53 + -87.4 = -140.4
	(b"11000010101001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011111001100110011010", b"11000011001010101100110011001101"), -- -83 + -87.8 = -170.8
	(b"11000000010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111111011001100110011010", b"11000010000011000110011001100111"), -- -3.4 + -31.7 = -35.1
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000101001100110011001101", b"11000010001101110011001100110100"), -- -8.6 + -37.2 = -45.8
	(b"01000010100000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001110111001100110011010", b"01000010111000010110011001100111"), -- 65.8 + 46.9 = 112.7
	(b"01000010100001110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110000011001100110011010", b"01000010101101111100110011001100"), -- 67.7 + 24.2 = 91.9
	(b"11000001000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110111001100110011010", b"11000010101011100011001100110100"), -- -9.3 + -77.8 = -87.1
	(b"11000010001000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011111001100110011010", b"11000011000000000110011001100110"), -- -40.6 + -87.8 = -128.4
	(b"01000010000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010001101100110011001101", b"11000001100000001100110011001110"), -- 33.6 + -49.7 = -16.1
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101011001100110011010", b"11000010101111111001100110011010"), -- -5 + -90.8 = -95.8
	(b"01000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101111010110011001100110", b"11000010101011100110011001100110"), -- 7.5 + -94.7 = -87.2
	(b"01000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100111100000000000000000", b"01000010101010000011001100110011"), -- 5.1 + 79 = 84.1
	(b"01000010011010111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110000100011001100110011", b"01000011000111000000000000000000"), -- 58.9 + 97.1 = 156
	(b"11000010101000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010001010011001100110011", b"11000011000000101000000000000000"), -- -81.2 + -49.3 = -130.5
	(b"11000010110000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001111000000000000000000", b"11000011000011111001100110011010"), -- -96.6 + -47 = -143.6
	(b"11000010100001010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101001010110011001100110", b"11000011000101010011001100110011"), -- -66.5 + -82.7 = -149.2
	(b"01000010010110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101000110000000000000000", b"11000001110111000000000000000000"), -- 54 + -81.5 = -27.5
	(b"01000010001001111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110001001100110011010", b"11000010010010011001100110011010"), -- 41.9 + -92.3 = -50.4
	(b"01000010001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111000000000000000000000", b"01000010100011100110011001100110"), -- 43.2 + 28 = 71.2
	(b"11000010101000100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101100100011001100110011", b"01000001000000000000000000000000"), -- -81.1 + 89.1 = 8
	(b"11000010101000001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010110001111001100110011010", b"11000011001101000001100110011010"), -- -80.3 + -99.8 = -180.1
	(b"01000010110001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001011011001100110011001101", b"01000010101001111001100110011001"), -- 98.6 + -14.8 = 83.8
	(b"10111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"11000000111100110011001100110011"), -- -0.9 + -6.7 = -7.6
	(b"01000001010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101101110011001100110011", b"01000010000100000110011001100110"), -- 13.2 + 22.9 = 36.1
	(b"01000010110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010011100000000000000000", b"01000011000100111000000000000000"), -- 96 + 51.5 = 147.5
	(b"01000010000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100010110011001100110011", b"11000010000100110011001100110011"), -- 32.8 + -69.6 = -36.8
	(b"11000010101111001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010010000000000000000", b"11000011001000101100110011001101"), -- -94.3 + -68.5 = -162.8
	(b"11000010010110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010010010011001100110011", b"11000010110100010011001100110011"), -- -54.3 + -50.3 = -104.6
	(b"01000010001011000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001100011001100110011", b"11000010011000000000000000000000"), -- 43.1 + -99.1 = -56
	(b"11000010100111010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011010110011001100110", b"11000011000101010110011001100110"), -- -78.7 + -70.7 = -149.4
	(b"11000010011000010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111001001100110011001101", b"11000001110111011001100110011001"), -- -56.3 + 28.6 = -27.7
	(b"11000010001001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101110000110011001100110", b"01000010010010111111111111111111"), -- -41.2 + 92.2 = 51
	(b"01000010011101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101010001100110011001101", b"01000010001000010011001100110100"), -- 61.4 + -21.1 = 40.3
	(b"01000010101011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001001010011001100110011", b"01000010001110100000000000000001"), -- 87.8 + -41.3 = 46.5
	(b"01000010100010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100000011001100110011", b"11000000001000000000000000000000"), -- 69.6 + -72.1 = -2.5
	(b"01000010000100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100001100000000000000000", b"01000010110011101100110011001101"), -- 36.4 + 67 = 103.4
	(b"11000010100111011100110011001101", b"00000000000000000000000000000000"),
	(b"10111101110011001100110011001101", b"11000010100111100000000000000000"), -- -78.9 + -0.1 = -79
	(b"01000010101000111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101110101100110011001101", b"11000001001110000000000000000000"), -- 81.9 + -93.4 = -11.5
	(b"01000010100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011011000000000000000000", b"01000011000001100011001100110011"), -- 75.2 + 59 = 134.2
	(b"11000001011101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010011101100110011001101", b"11000010100001100011001100110011"), -- -15.4 + -51.7 = -67.1
	(b"11000010100100110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001110100110011001100110", b"11000010111100001001100110011001"), -- -73.7 + -46.6 = -120.3
	(b"11000010110000011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110101000000000000000000", b"11000010111101101100110011001101"), -- -96.9 + -26.5 = -123.4
	(b"01000010101010000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010110000011100110011001101", b"01000011001101010000000000000000"), -- 84.1 + 96.9 = 181
	(b"11000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000001011011001100110011001101"), -- -5.3 + -9.5 = -14.8
	(b"01000010011110010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111001000000000000000000", b"01000010101101011001100110011010"), -- 62.3 + 28.5 = 90.8
	(b"11000010001010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101111111001100110011010", b"01000010010101100000000000000001"), -- -42.3 + 95.8 = 53.5
	(b"11000010101101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001011000011001100110011010", b"11000010100110011100110011001101"), -- -91 + 14.1 = -76.9
	(b"01000001011000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101101111100110011001101", b"01000010110101000000000000000000"), -- 14.1 + 91.9 = 106
	(b"11000001010101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001110100110011001100110", b"01000010000001010011001100110011"), -- -13.3 + 46.6 = 33.3
	(b"11000000011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010101000000000000000000", b"11000010011000111001100110011010"), -- -3.9 + -53 = -56.9
	(b"11000001101101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010110000010000000000000000", b"11000010111011101100110011001101"), -- -22.9 + -96.5 = -119.4
	(b"01000010110001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"01000010101111010011001100110011"), -- 98.2 + -3.6 = 94.6
	(b"01000010101101100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001101100110011001100110", b"01000010001101100000000000000000"), -- 91.1 + -45.6 = 45.5
	(b"01000001110110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"01000010000011100000000000000000"), -- 27.4 + 8.1 = 35.5
	(b"11000010110000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100100100011001100110011", b"11000001110000110011001100110100"), -- -97.5 + 73.1 = -24.4
	(b"01000001110111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100001100011001100110011", b"11000010000111011001100110011001"), -- 27.7 + -67.1 = -39.4
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111101001100110011001101", b"01000001110101001100110011001101"), -- -4 + 30.6 = 26.6
	(b"11000010100001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100011000000000000000000", b"11000011000010000000000000000000"), -- -66 + -70 = -136
	(b"01000010000100100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011001100110011001101", b"11000010010001111001100110011010"), -- 36.5 + -86.4 = -49.9
	(b"11000010011010000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001010011100110011001100110", b"11000010001101001100110011001100"), -- -58.1 + 12.9 = -45.2
	(b"11000001011010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100000100000000000000000", b"01000010010010010011001100110011"), -- -14.7 + 65 = 50.3
	(b"11000010100111010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110100110011001100110", b"10111111101100110011001101000000"), -- -78.6 + 77.2 = -1.4
	(b"01000010110001110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100111110110011001100110", b"01000011001100110110011001100110"), -- 99.7 + 79.7 = 179.4
	(b"11000001111000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100101011100110011001101", b"11000010110011100000000000000000"), -- -28.1 + -74.9 = -103
	(b"01000010000001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011000000000000000000", b"11000010010101000000000000000000"), -- 33 + -86 = -53
	(b"11000001000100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000011001100110011010", b"11000010110100111001100110011010"), -- -9 + -96.8 = -105.8
	(b"01000010100001000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101101111100110011001101", b"01000011000111100000000000000000"), -- 66.1 + 91.9 = 158
	(b"01000010001110010011001100110011", b"00000000000000000000000000000000"),
	(b"10111111111100110011001100110011", b"01000010001100011001100110011001"), -- 46.3 + -1.9 = 44.4
	(b"01000010000111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010000001100110011001101", b"01000010101011101100110011001101"), -- 39.2 + 48.2 = 87.4
	(b"11000010011110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000000100110011001100110", b"11000001111011001100110011001110"), -- -62.2 + 32.6 = -29.6
	(b"11000001101010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000111111001100110011010", b"01000001100101001100110011001110"), -- -21.3 + 39.9 = 18.6
	(b"01000010011011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101001100000000000000000", b"11000001101110110011001100110100"), -- 59.6 + -83 = -23.4
	(b"01000010100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011010000110011001100110", b"01000001100011110011001100110100"), -- 76 + -58.1 = 17.9
	(b"01000010000000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101110000011001100110011", b"01000010111110000110011001100110"), -- 32.1 + 92.1 = 124.2
	(b"01000001111010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111100000000000000000", b"11000010100000111001100110011010"), -- 29.2 + -95 = -65.8
	(b"11000010011010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"11000010100000001001100110011010"), -- -58.9 + -5.4 = -64.3
	(b"11000001011011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100111110011001100110011", b"11000010000010110011001100110011"), -- -14.9 + -19.9 = -34.8
	(b"11000010101100001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101111100110011001101", b"11000011001101000011001100110100"), -- -88.3 + -91.9 = -180.2
	(b"11000010100000010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010110000010000000000000000", b"01000010000000000000000000000000"), -- -64.5 + 96.5 = 32
	(b"11000010010001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"11000010001110110011001100110011"), -- -49.1 + 2.3 = -46.8
	(b"01000010100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011010100000000000000000", b"01000001001001001100110011010000"), -- 68.8 + -58.5 = 10.3
	(b"11000001100010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100101000000000000000000", b"11000010000011110011001100110011"), -- -17.3 + -18.5 = -35.8
	(b"11000010100101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100010100110011001100110", b"11000000100110011001100110100000"), -- -74 + 69.2 = -4.8
	(b"01000010010110111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010001001100110011010", b"01000011000010110011001100110100"), -- 54.9 + 84.3 = 139.2
	(b"11000010011001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010110001010011001100110011", b"01000010001001000110011001100110"), -- -57.5 + 98.6 = 41.1
	(b"01000010011001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111110001100110011001101", b"01000010101100010011001100110011"), -- 57.5 + 31.1 = 88.6
	(b"01000010001001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001010101100110011001100110", b"01000001110111110011001100110011"), -- 41.3 + -13.4 = 27.9
	(b"01000001101011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000100011001100110011010", b"01000010011010000110011001100111"), -- 21.7 + 36.4 = 58.1
	(b"01000010011110100000000000000000", b"00000000000000000000000000000000"),
	(b"11000000100000110011001100110011", b"01000010011010011001100110011010"), -- 62.5 + -4.1 = 58.4
	(b"11000010100101010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101000010110011001100110", b"01000000110000110011001100110000"), -- -74.6 + 80.7 = 6.1
	(b"01000010000100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001101000000000000000000", b"01000010101000110000000000000000"), -- 36.5 + 45 = 81.5
	(b"11000010000000100000000000000000", b"00000000000000000000000000000000"),
	(b"11000000001001100110011001100110", b"11000010000011000110011001100110"), -- -32.5 + -2.6 = -35.1
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001011001100110011001101", b"01000010001011000110011001100111"), -- -0.1 + 43.2 = 43.1
	(b"01000010101101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000010111001100110011010", b"01000010010111111001100110011010"), -- 90.8 + -34.9 = 55.9
	(b"11000010100111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001101111001100110011010", b"11000010111110110000000000000000"), -- -79.6 + -45.9 = -125.5
	(b"11000010100100000000000000000000", b"00000000000000000000000000000000"),
	(b"00111110100110011001100110011010", b"11000010100011110110011001100110"), -- -72 + 0.3 = -71.7
	(b"01000010001011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000010011001100110011", b"01000011000011000011001100110011"), -- 43.6 + 96.6 = 140.2
	(b"11000010100110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101010110000000000000000", b"11000011001000011110011001100110"), -- -76.4 + -85.5 = -161.9
	(b"11000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100101010110011001100110", b"11000010101000101001100110011001"), -- -6.6 + -74.7 = -81.3
	(b"01000010101010000011001100110011", b"00000000000000000000000000000000"),
	(b"01000001001110011001100110011010", b"01000010101111110110011001100110"), -- 84.1 + 11.6 = 95.7
	(b"01000010000011010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011011010011001100110011", b"01000010101111010011001100110011"), -- 35.3 + 59.3 = 94.6
	(b"11000010010010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010101001100110011010", b"01000001100110000000000000000010"), -- -50.3 + 69.3 = 19
	(b"11000010110001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111110011001100110011010", b"11000010100001111001100110011010"), -- -99 + 31.2 = -67.8
	(b"01000010000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000010000111011001100110011010"), -- 37.2 + 2.2 = 39.4
	(b"11000010100010101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010101100000000000000000", b"11000001011111001100110011010000"), -- -69.3 + 53.5 = -15.8
	(b"01000010101111101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111010100110011001100110", b"01000010111110010110011001100110"), -- 95.4 + 29.3 = 124.7
	(b"01000010101101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110110000000000000000", b"11000000001011001100110011000000"), -- 90.8 + -93.5 = -2.7
	(b"11000010101100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100110011001100110011010", b"11000010100011010011001100110100"), -- -89.8 + 19.2 = -70.6
	(b"11000010101101010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011100110011001100110", b"11000011001000011110011001100110"), -- -90.7 + -71.2 = -161.9
	(b"11000010101111111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010110001011100110011001101", b"11000011010000101011001100110100"), -- -95.8 + -98.9 = -194.7
	(b"01000010101110111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110000011100110011001101", b"01000011001111101011001100110100"), -- 93.8 + 96.9 = 190.7
	(b"01000010100100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101110110000000000000000", b"01000011001001101011001100110011"), -- 73.2 + 93.5 = 166.7
	(b"01000010011000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011100000000000000000", b"01000011000011110011001100110011"), -- 56.2 + 87 = 143.2
	(b"01000001111011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100011111001100110011010", b"01000010110010101001100110011010"), -- 29.5 + 71.8 = 101.3
	(b"11000001101001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011000101100110011001101", b"11000010100110110011001100110011"), -- -20.9 + -56.7 = -77.6
	(b"01000010010110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111000000000000000000000", b"01000010001111100110011001100110"), -- 54.6 + -7 = 47.6
	(b"11000010011010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011111000110011001100110", b"11000010111100101001100110011010"), -- -58.2 + -63.1 = -121.3
	(b"11000001101000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"11000001011001001100110011001110"), -- -20.2 + 5.9 = -14.3
	(b"01000010101011100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010110101100110011001101", b"01000010000000011001100110011001"), -- 87.1 + -54.7 = 32.4
	(b"11000010011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001010010011001100110011010", b"11000010100100101100110011001101"), -- -60.8 + -12.6 = -73.4
	(b"11000010011100010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110101001100110011001101", b"11000010101011011100110011001101"), -- -60.3 + -26.6 = -86.9
	(b"01000010101110101001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110100100110011001100110", b"01000010100001100000000000000000"), -- 93.3 + -26.3 = 67
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100011101001100110011010", b"01000010100110110110011001100111"), -- 6.4 + 71.3 = 77.7
	(b"11000010000011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101100001100110011001101", b"11000001010011100110011001100110"), -- -35 + 22.1 = -12.9
	(b"11000001101111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000011110011001100110011010", b"11000001110111100110011001100110"), -- -23.9 + -3.9 = -27.8
	(b"01000010101110010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010110000111100110011001101", b"01000011001111101000000000000000"), -- 92.6 + 97.9 = 190.5
	(b"11000010011010000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101111100110011001100110", b"01000010000101000110011001100110"), -- -58.1 + 95.2 = 37.1
	(b"11000001011111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001001110110011001100110011", b"11000000100001100110011001100110"), -- -15.9 + 11.7 = -4.2
	(b"01000010100110010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010100001100110011001101", b"01000011000000001110011001100110"), -- 76.7 + 52.2 = 128.9
	(b"11000010100101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011010100110011001100110", b"11000011000001100011001100110011"), -- -75.6 + -58.6 = -134.2
	(b"11000001110101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001100110001100110011001101", b"11000010001110000000000000000000"), -- -26.9 + -19.1 = -46
	(b"01000010001010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000001001100110011001101", b"01000010100110000000000000000000"), -- 42.8 + 33.2 = 76
	(b"01000010101000001001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101101100110011001100110", b"01000010011001100000000000000001"), -- 80.3 + -22.8 = 57.5
	(b"01000010010101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011011110011001100110011", b"11000000110010011001100110011000"), -- 53.5 + -59.8 = -6.3
	(b"11000010110000001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100100010000000000000000", b"11000001101111100110011001101000"), -- -96.3 + 72.5 = -23.8
	(b"01000001101101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011100001100110011001101", b"01000010101001100011001100110011"), -- 22.9 + 60.2 = 83.1
	(b"11000010100001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110000001100110011001101", b"11000010001011100000000000000000"), -- -67.6 + 24.1 = -43.5
	(b"01000001010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101011100011001100110011", b"11000010100100110000000000000000"), -- 13.6 + -87.1 = -73.5
	(b"01000001001010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001010110011001100110011010", b"01000001110000011001100110011010"), -- 10.6 + 13.6 = 24.2
	(b"01000001111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111110001100110011001101", b"01000010011011100000000000000000"), -- 28.4 + 31.1 = 59.5
	(b"11000001010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001111111100110011001100110", b"11000010001101000000000000000000"), -- -13.2 + -31.8 = -45
	(b"01000001110111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010101111001100110011010", b"11000001110100011001100110011010"), -- 27.7 + -53.9 = -26.2
	(b"11000001110110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100010101001100110011010", b"11000010110000010110011001100111"), -- -27.4 + -69.3 = -96.7
	(b"11000010100010101001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011001100110011001100110", b"11000010100100011100110011001101"), -- -69.3 + -3.6 = -72.9
	(b"01000010011010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101111110110011001100110", b"11000010000100111001100110011001"), -- 58.8 + -95.7 = -36.9
	(b"11000010100100001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001101000110011001100110", b"11000001110110011001100110011100"), -- -72.3 + 45.1 = -27.2
	(b"11000010100100010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100010110000000000000000", b"11000011000011100001100110011010"), -- -72.6 + -69.5 = -142.1
	(b"01000010011010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101110100110011001100110", b"11000010000010100110011001100110"), -- 58.6 + -93.2 = -34.6
	(b"01000010101110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011111111001100110011010", b"01000011000111000100110011001101"), -- 92.4 + 63.9 = 156.3
	(b"01000010101100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"01000010101111010011001100110100"), -- 89.8 + 4.8 = 94.6
	(b"01000010001000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101110000011001100110011", b"01000011000001010000000000000000"), -- 40.9 + 92.1 = 133
	(b"11000010101111000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001100001110011001100110011", b"11000010100110101001100110011001"), -- -94.2 + 16.9 = -77.3
	(b"11000010010001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001010110011001100110011010", b"11000010011110101100110011001100"), -- -49.1 + -13.6 = -62.7
	(b"01000010001011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"01000010001100011001100110011010"), -- 43.2 + 1.2 = 44.4
	(b"01000010010010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001111011001100110011010", b"01000000001001100110011001100000"), -- 50 + -47.4 = 2.6
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000000000000000000000", b"11000010100100110110011001100110"), -- 6.3 + -80 = -73.7
	(b"11000010101100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"11000010100111110000000000000000"), -- -89 + 9.5 = -79.5
	(b"01000010110001001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100111001001100110011010", b"01000011001100001001100110011010"), -- 98.3 + 78.3 = 176.6
	(b"11000001010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110111001100110011010", b"11000010110101101100110011001101"), -- -13.6 + -93.8 = -107.4
	(b"11000010101000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110100110011001100110", b"11000011001011100000000000000000"), -- -80.8 + -93.2 = -174
	(b"01000010101110010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111010001100110011001101", b"01000010011111100110011001100110"), -- 92.7 + -29.1 = 63.6
	(b"11000001001011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000111011001100110011010", b"01000001111001000000000000000001"), -- -10.9 + 39.4 = 28.5
	(b"11000010101001010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110111110011001100110011", b"11000010110111010011001100110011"), -- -82.7 + -27.9 = -110.6
	(b"11000010110001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010110011001100110011010", b"11000010001011100110011001100110"), -- -98 + 54.4 = -43.6
	(b"11000001110001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011011001100110011001101", b"01000010000010100110011001100110"), -- -24.6 + 59.2 = 34.6
	(b"11000010000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101001100110011001101", b"01000010010110110011001100110100"), -- -35.6 + 90.4 = 54.8
	(b"01000010100011000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011000111001100110011010", b"01000001010100011001100110011000"), -- 70 + -56.9 = 13.1
	(b"01000010010111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100010001001100110011010", b"01000010111101110000000000000000"), -- 55.2 + 68.3 = 123.5
	(b"01000010001100000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100001001001100110011010", b"01000010110111001100110011001101"), -- 44.1 + 66.3 = 110.4
	(b"11000001100110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010100000000000000000", b"01000010010001100110011001100110"), -- -19.4 + 69 = 49.6
	(b"11000010110001110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000011100110011001100110", b"11000011000001110001100110011010"), -- -99.5 + -35.6 = -135.1
	(b"01000010001011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011000101100110011001101", b"11000001010101001100110011001100"), -- 43.4 + -56.7 = -13.3
	(b"01000001101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110010100110011001100110", b"11000000011011001100110011001000"), -- 21.6 + -25.3 = -3.7
	(b"11000010000110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100010100000000000000000", b"01000001111100110011001100110100"), -- -38.6 + 69 = 30.4
	(b"01000010010100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001100010011001100110011010", b"01000010000011001100110011001101"), -- 52.4 + -17.2 = 35.2
	(b"01000010011001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101100000110011001100110", b"11000001111100111111111111111110"), -- 57.7 + -88.2 = -30.5
	(b"11000010110001000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011000100000000000000000", b"11000011000110101001100110011010"), -- -98.1 + -56.5 = -154.6
	(b"01000001110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101101000011001100110011", b"01000010111010000011001100110011"), -- 26 + 90.1 = 116.1
	(b"11000010000111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000001101100110011001101", b"11000010100100101100110011001101"), -- -39.7 + -33.7 = -73.4
	(b"11000010101111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100010000110011001100110", b"11000011001000111001100110011010"), -- -95.4 + -68.2 = -163.6
	(b"01000001100101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010101111001100110011010", b"11000010000011001100110011001101"), -- 18.7 + -53.9 = -35.2
	(b"11000010100100010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010010010011001100110011", b"11000001101100011001100110011010"), -- -72.5 + 50.3 = -22.2
	(b"01000001111110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010010000000000000000", b"01000010110001111100110011001101"), -- 31.4 + 68.5 = 99.9
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011100001100110011001101", b"01000010011111001100110011001101"), -- 3 + 60.2 = 63.2
	(b"01000010110001101001100110011010", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"01000010110001111100110011001101"), -- 99.3 + 0.6 = 99.9
	(b"01000001100001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101001010011001100110011", b"11000010100000110110011001100110"), -- 16.9 + -82.6 = -65.7
	(b"01000010101010000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100101101001100110011010", b"01000001000011001100110011001000"), -- 84.1 + -75.3 = 8.8
	(b"01000010100100101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001010000110011001100110011", b"01000010011101001100110011001101"), -- 73.4 + -12.2 = 61.2
	(b"01000010101100000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110010000000000000000", b"01000001001110011001100110011000"), -- 88.1 + -76.5 = 11.6
	(b"11000010000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100010110000000000000000", b"11000010110100100011001100110011"), -- -35.6 + -69.5 = -105.1
	(b"01000010110000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110000011001100110011010", b"01000010100100110011001100110100"), -- 97.8 + -24.2 = 73.6
	(b"11000001100010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001010001100110011001101", b"01000001110001100110011001100111"), -- -17.4 + 42.2 = 24.8
	(b"11000010101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011111100110011001100110", b"11000011000011111001100110011010"), -- -80 + -63.6 = -143.6
	(b"01000010100001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001010011001100110011", b"01000011000001010011001100110011"), -- 66.6 + 66.6 = 133.2
	(b"01000010100111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000000100110011001100110011", b"01000010100101110110011001100110"), -- 78 + -2.3 = 75.7
	(b"01000010110000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"01000010110101000000000000000000"), -- 97.8 + 8.2 = 106
	(b"01000001101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100100000011001100110011", b"01000010101110101001100110011010"), -- 21.2 + 72.1 = 93.3
	(b"01000010101111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110000110011001100110", b"01000001100110011001100110011100"), -- 95.4 + -76.2 = 19.2
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000000110011001100110", b"01000010100100001100110011001100"), -- -7.8 + 80.2 = 72.4
	(b"11000001100001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001100001100110011001100110", b"11000010000001101100110011001100"), -- -16.9 + -16.8 = -33.7
	(b"01000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101110010011001100110011", b"11000010101011100110011001100110"), -- 5.4 + -92.6 = -87.2
	(b"01000010001001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110001110011001100110011", b"01000001100001001100110011001101"), -- 41.5 + -24.9 = 16.6
	(b"11000010000011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100001001001100110011010", b"01000001111110011001100110011100"), -- -35.1 + 66.3 = 31.2
	(b"11000010110000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001010110000000000000000000", b"11000010101001011100110011001101"), -- -96.4 + 13.5 = -82.9
	(b"11000001001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000001100000011001100110011010"), -- -10.4 + -5.8 = -16.2
	(b"01000001111100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001001011100110011001100110", b"01000001100110011001100110011010"), -- 30.1 + -10.9 = 19.2
	(b"01000010001011101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000100110011001100110011", b"01000000110111001100110011010000"), -- 43.7 + -36.8 = 6.9
	(b"11000010011000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001010001100110011001100110", b"11000010001100011001100110011010"), -- -56.8 + 12.4 = -44.4
	(b"01000010000111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100101011100110011001101", b"01000010111001001100110011001101"), -- 39.5 + 74.9 = 114.4
	(b"11000010101101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010010110011001100110011", b"11000010000111001100110011001101"), -- -90 + 50.8 = -39.2
	(b"11000001111011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"11000010000111011001100110011010"), -- -29.9 + -9.5 = -39.4
	(b"01000010110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011101000110011001100110", b"01000011000111101011001100110011"), -- 97.6 + 61.1 = 158.7
	(b"01000001101001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101001010110011001100110", b"11000010011101110011001100110010"), -- 20.9 + -82.7 = -61.8
	(b"01000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110000110011001100110011", b"01000010111010101100110011001101"), -- 93 + 24.4 = 117.4
	(b"01000010101111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111011110011001100110011", b"01000010100000011100110011001101"), -- 94.8 + -29.9 = 64.9
	(b"01000010100111010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111001100110011001100110", b"01000010010001101100110011001101"), -- 78.5 + -28.8 = 49.7
	(b"01000010101101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110111001100110011010", b"11000000010000000000000000000000"), -- 90.8 + -93.8 = -3
	(b"01000010100110111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110000111001100110011010", b"01000011001011111001100110011010"), -- 77.8 + 97.8 = 175.6
	(b"01000010101001010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001101111001100110011010", b"01000011000000000110011001100110"), -- 82.5 + 45.9 = 128.4
	(b"01000010100000101100110011001101", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"01000010100000000011001100110011"), -- 65.4 + -1.3 = 64.1
	(b"11000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011110011001100110011010", b"11000010100010011100110011001101"), -- -6.5 + -62.4 = -68.9
	(b"01000010101101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001111001100110011001101", b"01000011000010100011001100110011"), -- 91 + 47.2 = 138.2
	(b"11000010011101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100101000110011001100110", b"01000001010011001100110011001000"), -- -61.4 + 74.2 = 12.8
	(b"01000001001010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100101001001100110011010", b"01000010101010011100110011001101"), -- 10.6 + 74.3 = 84.9
	(b"11000010100100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101100110011001100110011", b"11000010100001101100110011001101"), -- -73 + 5.6 = -67.4
	(b"01000010000010111001100110011010", b"00000000000000000000000000000000"),
	(b"01000000011011001100110011001101", b"01000010000110100110011001100111"), -- 34.9 + 3.7 = 38.6
	(b"01000010001110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010101100000000000000000", b"01000010110001111100110011001101"), -- 46.4 + 53.5 = 99.9
	(b"11000010101100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110001110011001100110011", b"11000011001110111001100110011010"), -- -88 + -99.6 = -187.6
	(b"01000010010001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011011100110011001101", b"01000011000010000001100110011010"), -- 49.2 + 86.9 = 136.1
	(b"01000010001000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100011110110011001100110", b"11000001111110110011001100110010"), -- 40.3 + -71.7 = -31.4
	(b"01000001111101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101000001100110011001101", b"01000010110111100110011001100110"), -- 30.8 + 80.4 = 111.2
	(b"01000010101101010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010110010011001100110011", b"01000010000100011001100110011001"), -- 90.7 + -54.3 = 36.4
	(b"01000010000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011001000110011001100110", b"11000001101100100110011001100110"), -- 34.8 + -57.1 = -22.3
	(b"01000010100000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011110100110011001100110", b"01000000001100110011001101000000"), -- 65.4 + -62.6 = 2.8
	(b"01000001111010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101100101001100110011010", b"01000010111011010110011001100111"), -- 29.4 + 89.3 = 118.7
	(b"01000010000101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101001011001100110011010", b"01000001100010011001100110011010"), -- 37.9 + -20.7 = 17.2
	(b"11000010110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100011001100110011001101", b"11000011001010000000000000000000"), -- -97.6 + -70.4 = -168
	(b"11000010100001000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010100101100110011001101", b"11000010111011011001100110011010"), -- -66.1 + -52.7 = -118.8
	(b"01000010101100001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100110111001100110011010", b"01000011001001100001100110011010"), -- 88.3 + 77.8 = 166.1
	(b"11000001101011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001001000000000000000000", b"11000010011110101100110011001101"), -- -21.7 + -41 = -62.7
	(b"01000010000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011100011001100110011010", b"01000010101111000000000000000000"), -- 33.6 + 60.4 = 94
	(b"11000010101111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000110101100110011001101", b"11000011000001001011001100110011"), -- -94 + -38.7 = -132.7
	(b"01000010100100010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001010001100110011001100110", b"01000010011100010011001100110010"), -- 72.7 + -12.4 = 60.3
	(b"01000001110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101010011001100110011", b"01000010100011011100110011001101"), -- 25.6 + 45.3 = 70.9
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101100110011001100110", b"01000010000101010011001100110011"), -- -8.3 + 45.6 = 37.3
	(b"11000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010011000000000000000000", b"01000010001010100110011001100110"), -- -8.4 + 51 = 42.6
	(b"01000001001111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100111100000000000000000", b"11000010100001100110011001100110"), -- 11.8 + -79 = -67.2
	(b"01000001101001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011100001100110011001101", b"11000010000111010011001100110100"), -- 20.9 + -60.2 = -39.3
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011000110011001100110011", b"01000010011010100110011001100110"), -- 1.8 + 56.8 = 58.6
	(b"11000001110001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101111011001100110011010", b"11000010111011110110011001100111"), -- -24.9 + -94.8 = -119.7
	(b"11000010001110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111110100110011001100110", b"11000010100110110000000000000000"), -- -46.2 + -31.3 = -77.5
	(b"11000010010110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001110011001100110011", b"01000001010101100110011001100100"), -- -54.2 + 67.6 = 13.4
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001010000000000000000000000", b"01000001010001100110011001100110"), -- 0.4 + 12 = 12.4
	(b"11000010101101001001100110011010", b"00000000000000000000000000000000"),
	(b"01000001001001001100110011001101", b"11000010101000000000000000000000"), -- -90.3 + 10.3 = -80
	(b"11000001110001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010110000010110011001100110", b"11000010111100101100110011001100"), -- -24.7 + -96.7 = -121.4
	(b"11000010101011001001100110011010", b"00000000000000000000000000000000"),
	(b"11000001011001001100110011001101", b"11000010110010010011001100110100"), -- -86.3 + -14.3 = -100.6
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001100000000000000000000", b"01000010000011101100110011001101"), -- -8.3 + 44 = 35.7
	(b"11000010100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101101100110011001101", b"01000001100000011001100110011100"), -- -75.2 + 91.4 = 16.2
	(b"11000001100110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111010110011001100110011", b"01000001001001100110011001100110"), -- -19 + 29.4 = 10.4
	(b"11000001100011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011001000000000000000000", b"01000010000111010011001100110011"), -- -17.7 + 57 = 39.3
	(b"01000010001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101110011100110011001101", b"11000010010100111001100110011010"), -- 40 + -92.9 = -52.9
	(b"11000001100010000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000001100001000000000000000000"), -- -17 + 0.5 = -16.5
	(b"11000010011001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011011111001100110011010", b"11000010111010100011001100110100"), -- -57.2 + -59.9 = -117.1
	(b"01000001110111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001100111001100110011010", b"11000001100010011001100110011010"), -- 27.7 + -44.9 = -17.2
	(b"01000010010010100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000001001100110011001101", b"01000010011010110011001100110011"), -- 50.5 + 8.3 = 58.8
	(b"11000010000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110001100110011001100110", b"11000010011110011001100110011001"), -- -37.6 + -24.8 = -62.4
	(b"01000001011100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010010100000000000000000", b"11000010000011011001100110011010"), -- 15.1 + -50.5 = -35.4
	(b"11000010001000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000111000110011001100110", b"10111111110110011001100110100000"), -- -40.8 + 39.1 = -1.7
	(b"11000010100100011100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000000110011001100110011", b"11000010100000010110011001100111"), -- -72.9 + 8.2 = -64.7
	(b"11000001011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101100011001100110011", b"11000010110101010110011001100110"), -- -15.6 + -91.1 = -106.7
	(b"11000010011001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101110100110011001100110", b"11000011000101110000000000000000"), -- -57.8 + -93.2 = -151
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110001110011001100110011", b"11000001100101100110011001100110"), -- 6.1 + -24.9 = -18.8
	(b"11000010010011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111011100110011001100110", b"11000001101011001100110011001110"), -- -51.4 + 29.8 = -21.6
	(b"11000010100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001001001100110011001101", b"11000010000000011001100110011001"), -- -73.6 + 41.2 = -32.4
	(b"11000010100100101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000010000110011001100110", b"11000010000111010011001100110100"), -- -73.4 + 34.1 = -39.3
	(b"01000010110000110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110001000000000000000000", b"01000011010000111011001100110011"), -- 97.7 + 98 = 195.7
	(b"01000010001010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100101100110011001100110", b"01000010000101111001100110011001"), -- 42.6 + -4.7 = 37.9
	(b"11000010011100101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101011011001100110011010", b"11000010000111000000000000000000"), -- -60.7 + 21.7 = -39
	(b"01000010100001110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100101001001100110011010", b"11000000110110011001100110100000"), -- 67.5 + -74.3 = -6.8
	(b"11000010000110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101111010000000000000000", b"01000010011000100000000000000000"), -- -38 + 94.5 = 56.5
	(b"11000010101110110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100011100110011001100110", b"11000001101101000000000000000000"), -- -93.7 + 71.2 = -22.5
	(b"11000001111111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001101100110011001100110", b"11000010100110110000000000000000"), -- -31.9 + -45.6 = -77.5
	(b"01000001101011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001001011001100110011010", b"11000001100111000000000000000001"), -- 21.9 + -41.4 = -19.5
	(b"01000010100100110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001001010110011001100110011", b"01000010101010001100110011001100"), -- 73.7 + 10.7 = 84.4
	(b"11000010000011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100101001100110011010", b"11000010110110100011001100110100"), -- -35.8 + -73.3 = -109.1
	(b"01000001001011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101111110011001100110011", b"11000010101010010110011001100110"), -- 10.9 + -95.6 = -84.7
	(b"01000010100111010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011011100110011001100110", b"01000001100110001100110011001100"), -- 78.7 + -59.6 = 19.1
	(b"01000001101101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001100000000000000000000", b"01000010100001011001100110011010"), -- 22.8 + 44 = 66.8
	(b"01000000110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111100110011001100110011", b"01000010000101010011001100110011"), -- 6.9 + 30.4 = 37.3
	(b"11000001101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011111100000000000000000", b"11000010101011001001100110011010"), -- -22.8 + -63.5 = -86.3
	(b"11000010101111100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111100110011001100110011", b"11000010111110101100110011001101"), -- -95 + -30.4 = -125.4
	(b"11000000000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001000111001100110011010", b"11000010001011010011001100110100"), -- -2.4 + -40.9 = -43.3
	(b"11000001011001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111011011001100110011010", b"01000001011101100110011001100111"), -- -14.3 + 29.7 = 15.4
	(b"01000001100010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110011001100110011001101", b"11000001000001001100110011001110"), -- 17.3 + -25.6 = -8.3
	(b"11000010101000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010000010011001100110011", b"11000011000000001110011001100110"), -- -80.6 + -48.3 = -128.9
	(b"11000010011011010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100101100110011001100110", b"11000011000001101000000000000000"), -- -59.3 + -75.2 = -134.5
	(b"11000010010101000110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100000000000000000000000", b"11000010010001000110011001100110"), -- -53.1 + 4 = -49.1
	(b"11000010001110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100000110011001100110011", b"11000001111100001100110011001101"), -- -46.5 + 16.4 = -30.1
	(b"11000001110111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101111001100110011010", b"01000010100000000000000000000000"), -- -27.8 + 91.8 = 64
	(b"01000010011100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100110010000000000000000", b"11000001100000110011001100110100"), -- 60.1 + -76.5 = -16.4
	(b"01000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011011100110011001101", b"11000010100000100110011001100111"), -- 5.7 + -70.9 = -65.2
	(b"01000010110001000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101100111100110011001101", b"01000001000000110011001100110000"), -- 98.1 + -89.9 = 8.2
	(b"11000001111101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001010101100110011001101", b"11000010100100110011001100110011"), -- -30.9 + -42.7 = -73.6
	(b"01000000110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010110001100110011001101", b"01000010011100101100110011001101"), -- 6.5 + 54.2 = 60.7
	(b"11000001010100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000101001100110011010", b"11000010101111001100110011001101"), -- -13.1 + -81.3 = -94.4
	(b"01000010010000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000000000000000000000000", b"01000010101000010110011001100110"), -- 48.7 + 32 = 80.7
	(b"01000001110001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101100010110011001100110", b"11000010100000000011001100110011"), -- 24.6 + -88.7 = -64.1
	(b"01000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011100000110011001100110", b"01000011000110010001100110011010"), -- 93 + 60.1 = 153.1
	(b"11000010100111011100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"11000010100111001100110011001101"), -- -78.9 + 0.5 = -78.4
	(b"01000010110000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110000100110011001100110", b"01000010100100100011001100110100"), -- 97.4 + -24.3 = 73.1
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010101110011001100110011", b"01000010001110010011001100110011"), -- -7.5 + 53.8 = 46.3
	(b"01000010100010111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101101010000000000000000", b"01000011001000000110011001100110"), -- 69.9 + 90.5 = 160.4
	(b"11000010010111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100010111100110011001101", b"11000010111110110000000000000000"), -- -55.6 + -69.9 = -125.5
	(b"01000010110000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001111110011001100110011", b"01000011000100000000000000000000"), -- 96.2 + 47.8 = 144
	(b"11000010101001011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101010111100110011001101", b"11000011001010001100110011001101"), -- -82.9 + -85.9 = -168.8
	(b"11000010101000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010001001100110011010", b"11000001010101001100110011001000"), -- -81.6 + 68.3 = -13.3
	(b"01000010000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000111011001100110011010", b"10111111111001100110011010000000"), -- 37.6 + -39.4 = -1.8
	(b"11000010000011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000010010011001100110011", b"10111111100011001100110011100000"), -- -35.4 + 34.3 = -1.1
	(b"01000010011010100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101111100110011001101", b"11000010000001011001100110011010"), -- 58.5 + -91.9 = -33.4
	(b"11000001010111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111111001100110011001101", b"11000000101111001100110011001101"), -- -13.8 + 7.9 = -5.9
	(b"01000001111001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000100101100110011001101", b"11000000111110011001100110011100"), -- 28.9 + -36.7 = -7.8
	(b"11000010000011111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001101101001100110011001101", b"11000001010101001100110011001110"), -- -35.9 + 22.6 = -13.3
	(b"11000010001101111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101100010110011001100110", b"01000010001010110011001100110010"), -- -45.9 + 88.7 = 42.8
	(b"01000010000101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010001001100110011010", b"11000010001110100000000000000001"), -- 37.8 + -84.3 = -46.5
	(b"11000001101000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111010011001100110011", b"01000010000011010011001100110011"), -- -20 + 55.3 = 35.3
	(b"01000010010111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111100000000000000000000", b"01000001110010001100110011001100"), -- 55.1 + -30 = 25.1
	(b"01000010011101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010011001100110011001101", b"01000010100000010110011001100110"), -- 61.5 + 3.2 = 64.7
	(b"11000010100100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000011100110011001100110", b"11000010110110100110011001100110"), -- -73.6 + -35.6 = -109.2
	(b"01000010100011110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101000000000000000000000", b"01000011000101111000000000000000"), -- 71.5 + 80 = 151.5
	(b"11000010101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100100000000000000000000", b"11000011001000110011001100110011"), -- -91.2 + -72 = -163.2
	(b"01000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001001000000000000000000", b"01000010001111010011001100110011"), -- 6.3 + 41 = 47.3
	(b"11000010001111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"11000010001101101100110011001101"), -- -47.8 + 2.1 = -45.7
	(b"11000010100100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000111000110011001100110", b"11000010110111101001100110011001"), -- -72.2 + -39.1 = -111.3
	(b"01000010101000010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011101001100110011010", b"11000000110110011001100110100000"), -- 80.5 + -87.3 = -6.8
	(b"01000010001011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001101101100110011001101", b"11000000000011001100110011010000"), -- 43.5 + -45.7 = -2.2
	(b"11000001101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100101100110011001100110", b"01000010010101111111111111111111"), -- -21.2 + 75.2 = 54
	(b"01000001101010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010110001100110011001101", b"11000010000001000110011001100110"), -- 21.1 + -54.2 = -33.1
	(b"11000001101100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101111000000000000000000", b"11000010001101110011001100110011"), -- -22.3 + -23.5 = -45.8
	(b"11000001010110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000111100110011001100110", b"11000010010101010011001100110011"), -- -13.7 + -39.6 = -53.3
	(b"01000001101001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001000111001100110011010", b"11000001101000011001100110011010"), -- 20.7 + -40.9 = -20.2
	(b"11000010101000001001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111000011001100110011010", b"11000010010100000110011001100111"), -- -80.3 + 28.2 = -52.1
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001011001100110011001100110", b"01000001011111100110011001100110"), -- 1.5 + 14.4 = 15.9
	(b"01000010000010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011001101100110011001101", b"01000010101110000000000000000000"), -- 34.3 + 57.7 = 92
	(b"01000001101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001001001100110011010", b"11000010100101110000000000000000"), -- 22.8 + -98.3 = -75.5
	(b"01000010110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010001100110011001100110", b"01000010010000000000000000000000"), -- 97.6 + -49.6 = 48
	(b"01000010010011100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100000100110011001100110", b"01000010100001111001100110011010"), -- 51.5 + 16.3 = 67.8
	(b"11000010010000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000001000000000000000000", b"11000010101000101100110011001101"), -- -48.4 + -33 = -81.4
	(b"01000010100000100011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101001011001100110011010", b"01000010001100011001100110011001"), -- 65.1 + -20.7 = 44.4
	(b"01000001110101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111001001100110011001101", b"01000010010111100000000000000000"), -- 26.9 + 28.6 = 55.5
	(b"11000010011101101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101011011001100110011010", b"11000010001000000000000000000000"), -- -61.7 + 21.7 = -40
	(b"11000010011010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001111110011001100110011010", b"11000001110110110011001100110010"), -- -58.6 + 31.2 = -27.4
	(b"01000010101000000011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101110110011001100110011", b"01000010011000101100110011001100"), -- 80.1 + -23.4 = 56.7
	(b"01000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101000000110011001100110", b"11000010100111000011001100110011"), -- 2.1 + -80.2 = -78.1
	(b"11000001110000100110011001100110", b"00000000000000000000000000000000"),
	(b"10111111111001100110011001100110", b"11000001110100001100110011001100"), -- -24.3 + -1.8 = -26.1
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010101001100110011001101", b"11000010011101111001100110011010"), -- -8.7 + -53.2 = -61.9
	(b"01000010001001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111100011001100110011010", b"01000010100100000011001100110100"), -- 41.9 + 30.2 = 72.1
	(b"11000001111010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000010110011001100110011", b"01000000101100000000000000000000"), -- -29.3 + 34.8 = 5.5
	(b"01000010101101110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011101000000000000000000", b"01000011000110001011001100110011"), -- 91.7 + 61 = 152.7
	(b"11000010101110010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000000011001100110011010", b"11000010101010001100110011001101"), -- -92.5 + 8.1 = -84.4
	(b"11000001100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101110100110011001100110", b"11000010001000100000000000000000"), -- -17.2 + -23.3 = -40.5
	(b"11000001100001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"11000001000100000000000000000000"), -- -16.5 + 7.5 = -9
	(b"01000010101000010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000010101100101001100110011010"), -- 80.5 + 8.8 = 89.3
	(b"11000010010101101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100100010110011001100110", b"11000010111111001100110011001100"), -- -53.7 + -72.7 = -126.4
	(b"01000010101000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000010101011110011001100110100"), -- 80.8 + 6.8 = 87.6
	(b"11000001101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100000010000000000000000", b"11000010101010011100110011001101"), -- -20.4 + -64.5 = -84.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011010101100110011001101", b"01000010011101100000000000000000"), -- 2.8 + 58.7 = 61.5
	(b"11000010000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101010111001100110011010", b"01000010010010001100110011001110"), -- -35.6 + 85.8 = 50.2
	(b"01000010110001000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011101100110011001100110", b"01000011000111111011001100110011"), -- 98.1 + 61.6 = 159.7
	(b"01000010011001011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101111110011001100110011", b"01000011000110010000000000000000"), -- 57.4 + 95.6 = 153
	(b"11000001100110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011101011001100110011010", b"01000010001010000110011001100111"), -- -19.3 + 61.4 = 42.1
	(b"11000010000111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111000110011001100110011", b"11000001001100000000000000000010"), -- -39.4 + 28.4 = -11
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011000100110011001100110", b"11000010100000101001100110011001"), -- -8.7 + -56.6 = -65.3
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110011110011001100110011", b"11000001100101000000000000000000"), -- 7.4 + -25.9 = -18.5
	(b"11000010101011000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101111010110011001100110", b"11000011001101001011001100110011"), -- -86 + -94.7 = -180.7
	(b"01000001110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111000000000000000000", b"01000010101000100000000000000000"), -- 26 + 55 = 81
	(b"11000010100110111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010111000000000000000000", b"11000001101101110011001100110100"), -- -77.9 + 55 = -22.9
	(b"11000001111100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011001000000000000000000", b"01000001110101110011001100110011"), -- -30.1 + 57 = 26.9
	(b"01000010011111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010000110011001100110", b"11000000100110011001100110010000"), -- 63.4 + -68.2 = -4.8
	(b"01000001110111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001011010011001100110011010", b"01000001010101001100110011001100"), -- 27.9 + -14.6 = 13.3
	(b"01000010101101010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101110001001100110011010", b"10111111110011001100110100000000"), -- 90.7 + -92.3 = -1.60001
	(b"01000010100010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001000000110011001100110", b"01000010110110011100110011001101"), -- 68.8 + 40.1 = 108.9
	(b"01000010101000001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001010100000000000000000", b"01000010000101110011001100110100"), -- 80.3 + -42.5 = 37.8
	(b"11000010011110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001010001100110011001101", b"11000010110100100011001100110100"), -- -62.9 + -42.2 = -105.1
	(b"11000010011000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010000100110011001100110", b"11000010110100110000000000000000"), -- -56.9 + -48.6 = -105.5
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110110100110011001100110", b"11000001111110000000000000000000"), -- -3.7 + -27.3 = -31
	(b"11000010011001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000100100000000000000000", b"11000010101111000000000000000000"), -- -57.5 + -36.5 = -94
	(b"01000010001011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001111000110011001100110", b"01000010101101000110011001100110"), -- 43.1 + 47.1 = 90.2
	(b"01000001111001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001100111001100110011010", b"01000010100100110000000000000000"), -- 28.6 + 44.9 = 73.5
	(b"11000001100001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000011111001100110011010", b"11000010010100100110011001100111"), -- -16.7 + -35.9 = -52.6
	(b"11000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110010001100110011001101", b"11000001111100000000000000000000"), -- -4.9 + -25.1 = -30
	(b"11000010011110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011001000110011001100110", b"11000010111011101100110011001100"), -- -62.3 + -57.1 = -119.4
	(b"11000001110011100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000001110100011001100110011001"), -- -25.8 + -0.4 = -26.2
	(b"01000010000010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"01000001110110001100110011001101"), -- 34.2 + -7.1 = 27.1
	(b"01000010001011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"01000010000010100000000000000000"), -- 43.5 + -9 = 34.5
	(b"01000010101111110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001110111001100110011010", b"01000010010000110011001100110010"), -- 95.7 + -46.9 = 48.8
	(b"11000010000010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100010110011001100110011", b"11000001100001100110011001100111"), -- -34.2 + 17.4 = -16.8
	(b"01000010000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001011001100110011001101", b"01000010000011100000000000000000"), -- 32.8 + 2.7 = 35.5
	(b"11000001111111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100001010000000000000000", b"11000010110001001100110011001101"), -- -31.9 + -66.5 = -98.4
	(b"11000010110000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101111000110011001100110", b"11000000011001100110011010000000"), -- -97.8 + 94.2 = -3.60001
	(b"01000010110000001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110001000011001100110011", b"01000011010000100110011001100110"), -- 96.3 + 98.1 = 194.4
	(b"01000010001110101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010110001000110011001100110", b"11000010010011011111111111111111"), -- 46.7 + -98.2 = -51.5
	(b"01000010100110011100110011001101", b"00000000000000000000000000000000"),
	(b"10111111100011001100110011001101", b"01000010100101111001100110011010"), -- 76.9 + -1.1 = 75.8
	(b"01000010001111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110100100110011001100110", b"01000001101001100110011001100110"), -- 47.1 + -26.3 = 20.8
	(b"01000010001100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001011011001100110011010", b"00111111001100110011001100000000"), -- 44.1 + -43.4 = 0.699997
	(b"01000010110001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101100011001100110011010", b"01000011001110101100110011001101"), -- 98 + 88.8 = 186.8
	(b"11000010101001100011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101101000000000000000000", b"11000010110100110011001100110011"), -- -83.1 + -22.5 = -105.6
	(b"11000010100010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001110100000000000000000", b"11000010111010001001100110011010"), -- -69.8 + -46.5 = -116.3
	(b"11000010101001110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110110011001100110011010", b"11000010110111011100110011001100"), -- -83.7 + -27.2 = -110.9
	(b"11000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000100101100110011001101", b"11000010001110001100110011001101"), -- -9.5 + -36.7 = -46.2
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"11000000110111111111111111111111"), -- -8.9 + 1.9 = -7
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000000100000000000000000", b"01000001111000110011001100110011"), -- -4.1 + 32.5 = 28.4
	(b"01000001111011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100100001001100110011010", b"01000010110011000110011001100111"), -- 29.9 + 72.3 = 102.2
	(b"01000010011000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000011001100110011001101", b"01000001101010110011001100110010"), -- 56.6 + -35.2 = 21.4
	(b"11000001111111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100010001100110011001101", b"01000010000100101100110011001101"), -- -31.7 + 68.4 = 36.7
	(b"11000001111101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001011001100110011001100110", b"11000001100000100110011001100111"), -- -30.7 + 14.4 = -16.3
	(b"01000010011101101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011010010011001100110011", b"01000010111100000000000000000000"), -- 61.7 + 58.3 = 120
	(b"11000001110100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100101001100110011001101", b"11000000111100000000000000000000"), -- -26.1 + 18.6 = -7.5
	(b"01000010110001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100010011001100110011010", b"01000001111100011001100110011000"), -- 99 + -68.8 = 30.2
	(b"01000010100111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000010001100110011001101", b"01000010111001000000000000000000"), -- 79.8 + 34.2 = 114
	(b"01000001101111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100001100011001100110011", b"11000010001011001100110011001100"), -- 23.9 + -67.1 = -43.2
	(b"11000010100101010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101010011001100110011", b"01000001011111100110011001101000"), -- -74.7 + 90.6 = 15.9
	(b"01000010001010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001011100011001100110011010", b"01000010011001101100110011001100"), -- 42.6 + 15.1 = 57.7
	(b"01000001101101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111000100110011001100110", b"01000010010011001100110011001100"), -- 22.9 + 28.3 = 51.2
	(b"01000010011011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000111100110011001101", b"01000011000111010000000000000000"), -- 59.1 + 97.9 = 157
	(b"01000010100100110000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111001100110011001100110", b"01000010110011001001100110011010"), -- 73.5 + 28.8 = 102.3
	(b"11000010101110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100001100110011001100110", b"11000010100110010011001100110100"), -- -93.4 + 16.8 = -76.6
	(b"11000001100001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110110110011001100110", b"01000010011100111001100110011001"), -- -16.8 + 77.7 = 60.9
	(b"01000010001010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"01000010000010011001100110011010"), -- 42.2 + -7.8 = 34.4
	(b"11000010001100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101110000000000000000000", b"11000011000010000011001100110011"), -- -44.2 + -92 = -136.2
	(b"01000001101010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000001111000110011001100110011"), -- 21.3 + 7.1 = 28.4
	(b"11000010101111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011001010011001100110011", b"11000011000110000001100110011010"), -- -94.8 + -57.3 = -152.1
	(b"01000010100110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010001001100110011010", b"01000001000110000000000000000000"), -- 77.8 + -68.3 = 9.5
	(b"01000010001011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001111100000000000000000", b"11000000011011001100110011010000"), -- 43.8 + -47.5 = -3.7
	(b"01000010011110000000000000000000", b"00000000000000000000000000000000"),
	(b"00111111001100110011001100110011", b"01000010011110101100110011001101"), -- 62 + 0.7 = 62.7
	(b"01000010101111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011100110011001100110", b"01000001101110000000000000000000"), -- 94.2 + -71.2 = 23
	(b"11000010010000100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100111110000000000000000", b"11000011000000000000000000000000"), -- -48.5 + -79.5 = -128
	(b"01000010011111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110001010000000000000000", b"01000011001000100110011001100110"), -- 63.9 + 98.5 = 162.4
	(b"01000010001110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110010000000000000000000", b"01000010100011110011001100110011"), -- 46.6 + 25 = 71.6
	(b"11000010100000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011101000110011001100110", b"11000010111111010000000000000000"), -- -65.4 + -61.1 = -126.5
	(b"11000001001010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010110111001100110011010", b"01000010001100001100110011001101"), -- -10.7 + 54.9 = 44.2
	(b"11000000011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010010010011001100110011", b"01000010001110100110011001100110"), -- -3.7 + 50.3 = 46.6
	(b"11000010001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010101001100110011001101", b"11000010110001000000000000000000"), -- -44.8 + -53.2 = -98
	(b"01000010000001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"01000001101110100110011001100110"), -- 33 + -9.7 = 23.3
	(b"11000010101100101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100000100011001100110011", b"11000011000110101000000000000000"), -- -89.4 + -65.1 = -154.5
	(b"11000010110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110100011001100110011010", b"11000010100010111001100110011010"), -- -96 + 26.2 = -69.8
	(b"01000010001111010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001010110110011001100110011", b"01000010000001100110011001100110"), -- 47.3 + -13.7 = 33.6
	(b"01000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000001010011001100110011", b"01000010000100110011001100110011"), -- 3.5 + 33.3 = 36.8
	(b"01000001110111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111111000000000000000000", b"01000010011011000000000000000000"), -- 27.5 + 31.5 = 59
	(b"11000010100111010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"11000010100010110110011001100110"), -- -78.5 + 8.8 = -69.7
	(b"11000010101101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000001001100110011001101", b"11000010110010000011001100110100"), -- -91.8 + -8.3 = -100.1
	(b"01000010011100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101111000011001100110011", b"01000011000110101001100110011010"), -- 60.5 + 94.1 = 154.6
	(b"01000010100101010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100101011001100110011010", b"01000011000101011000000000000000"), -- 74.7 + 74.8 = 149.5
	(b"11000010101111010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011000000000000000000", b"11000011001001001011001100110011"), -- -94.7 + -70 = -164.7
	(b"11000001110100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110001001100110011001101", b"11000010010010100110011001100110"), -- -26 + -24.6 = -50.6
	(b"11000010001110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000000000000000000000", b"01000010010001010011001100110011"), -- -46.7 + 96 = 49.3
	(b"01000010101110101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101110100000000000000000", b"00111110110011001100110100000000"), -- 93.4 + -93 = 0.400002
	(b"11000010010100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001000111001100110011010", b"11000010101110101001100110011010"), -- -52.4 + -40.9 = -93.3
	(b"01000010110001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100101011001100110011010", b"01000010111011000011001100110100"), -- 99.4 + 18.7 = 118.1
	(b"11000010101100101001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000101101100110011001101", b"11000010111111100000000000000000"), -- -89.3 + -37.7 = -127
	(b"10111111110110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001100100110011001100110", b"11000010001110010011001100110011"), -- -1.7 + -44.6 = -46.3
	(b"11000001111011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000101000110011001100110011", b"11000010000010110011001100110011"), -- -29.7 + -5.1 = -34.8
	(b"01000010011101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001001011001100110011010", b"01000001101000001100110011001100"), -- 61.5 + -41.4 = 20.1
	(b"11000010100111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011100110011001100110", b"11000011001001100110011001100110"), -- -79.2 + -87.2 = -166.4
	(b"11000010100000010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100101110000000000000000", b"01000001001011001100110011010000"), -- -64.7 + 75.5 = 10.8
	(b"11000000101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011000101100110011001101", b"11000010011101101100110011001101"), -- -5 + -56.7 = -61.7
	(b"01000010101101011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000011100110011001101", b"01000001001000000000000000000000"), -- 90.9 + -80.9 = 10
	(b"01000010100110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011111000110011001100110", b"01000001010110000000000000000000"), -- 76.6 + -63.1 = 13.5
	(b"11000001101100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010011101100110011001101", b"01000001111010110011001100110100"), -- -22.3 + 51.7 = 29.4
	(b"01000010100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101001100110011001101", b"11000001101110011001100110011100"), -- 67.2 + -90.4 = -23.2
	(b"11000010101001010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100111000011001100110011", b"11000000100011001100110011010000"), -- -82.5 + 78.1 = -4.4
	(b"11000010010110000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001100011000000000000000000", b"11000010000100100110011001100110"), -- -54.1 + 17.5 = -36.6
	(b"11000010101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100100000011001100110011", b"11000001010010110011001100111000"), -- -84.8 + 72.1 = -12.7
	(b"01000001001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101110110011001100110011", b"11000010101001001100110011001101"), -- 11.2 + -93.6 = -82.4
	(b"01000010001111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101101010110011001100110", b"01000011000010101001100110011010"), -- 47.9 + 90.7 = 138.6
	(b"11000001110000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100011000011001100110011", b"01000010001101111001100110011001"), -- -24.2 + 70.1 = 45.9
	(b"11000010010100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101000000000000000000000", b"11000010100100010011001100110011"), -- -52.6 + -20 = -72.6
	(b"11000010011001000110011001100110", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000010011001110011001100110011"), -- -57.1 + -0.7 = -57.8
	(b"11000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101011000000000000000000", b"01000001010011001100110011001101"), -- -8.7 + 21.5 = 12.8
	(b"11000010010011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100010000000000000000000", b"11000010000010101100110011001101"), -- -51.7 + 17 = -34.7
	(b"01000010110001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001111100000000000000000", b"01000011000100100001100110011010"), -- 98.6 + 47.5 = 146.1
	(b"01000000110101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011011100110011001100110", b"11000001000000110011001100110011"), -- 6.7 + -14.9 = -8.2
	(b"01000010100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100000000011001100110011", b"01000001011001001100110011010000"), -- 78.4 + -64.1 = 14.3
	(b"11000010001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000111110011001100110011", b"11000010100111111001100110011010"), -- -40 + -39.8 = -79.8
	(b"11000010100000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100100001100110011001101", b"01000000111000000000000000000000"), -- -65.4 + 72.4 = 7
	(b"11000010100000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000010100000000000000000", b"11000010110001010110011001100110"), -- -64.2 + -34.5 = -98.7
	(b"11000001010110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100000100011001100110011", b"01000010010011011001100110011001"), -- -13.7 + 65.1 = 51.4
	(b"01000010010111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011100011001100110011010", b"11000000101011001100110011010000"), -- 55 + -60.4 = -5.4
	(b"01000001011010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101101110000000000000000", b"01000010110101000000000000000000"), -- 14.5 + 91.5 = 106
	(b"01000010000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010011100110011001100110", b"01000010101010100110011001100110"), -- 33.6 + 51.6 = 85.2
	(b"01000010110001110011001100110011", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000010110010000000000000000000"), -- 99.6 + 0.4 = 100
	(b"01000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101100000000000000000000", b"01000010110000000110011001100110"), -- 8.2 + 88 = 96.2
	(b"01000010100001011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001011101100110011001100110", b"01000010010011100000000000000000"), -- 66.9 + -15.4 = 51.5
	(b"01000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100111000000000000000000", b"11000001010111001100110011001101"), -- 5.7 + -19.5 = -13.8
	(b"11000010001110101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111110001100110011001101", b"11000010100110111001100110011010"), -- -46.7 + -31.1 = -77.8
	(b"11000010000000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000110000000000000000000", b"01000000101110011001100110011000"), -- -32.2 + 38 = 5.8
	(b"01000010101100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010110010011001100110011", b"01000010000010000110011001100111"), -- 88.4 + -54.3 = 34.1
	(b"01000010011010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001010110000000000000000000", b"01000010001100111001100110011010"), -- 58.4 + -13.5 = 44.9
	(b"01000010100100010110011001100110", b"00000000000000000000000000000000"),
	(b"01000001010000000000000000000000", b"01000010101010010110011001100110"), -- 72.7 + 12 = 84.7
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001010001100110011001101", b"11000010000011110011001100110011"), -- 6.4 + -42.2 = -35.8
	(b"01000001100000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010010010011001100110011", b"11000010000010001100110011001100"), -- 16.1 + -50.3 = -34.2
	(b"01000010101101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101110001100110011001101", b"11000000000000000000000000000000"), -- 90.4 + -92.4 = -2
	(b"01000010011000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111010110011001100110011", b"01000010101011000011001100110011"), -- 56.7 + 29.4 = 86.1
	(b"11000010011011010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101000000000000000000", b"01000001011010110011001100110100"), -- -59.3 + 74 = 14.7
	(b"11000010011111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011011010011001100110011", b"11000000100100000000000000000000"), -- -63.8 + 59.3 = -4.5
	(b"11000001100010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010010001100110011001101", b"01000010000000110011001100110100"), -- -17.4 + 50.2 = 32.8
	(b"01000010001110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111000110011001100110011", b"01000010000111000110011001100111"), -- 46.2 + -7.1 = 39.1
	(b"01000010000000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101000000011001100110011", b"01000010111000011100110011001100"), -- 32.8 + 80.1 = 112.9
	(b"11000010101101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011011100110011001100110", b"11000011000101100000000000000000"), -- -90.4 + -59.6 = -150
	(b"11000001111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111110100110011001100110", b"11000010011100000110011001100110"), -- -28.8 + -31.3 = -60.1
	(b"01000010100100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110110000000000000000000", b"01000010110010000110011001100110"), -- 73.2 + 27 = 100.2
	(b"11000010001101000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000101011001100110011010", b"11000010101001010000000000000000"), -- -45.1 + -37.4 = -82.5
	(b"11000000101111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101110000110011001100110", b"01000010101011001001100110011001"), -- -5.9 + 92.2 = 86.3
	(b"01000010000001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010011111001100110011010", b"01000010101010111001100110011010"), -- 33.9 + 51.9 = 85.8
	(b"11000010100001111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000000110011001100110011", b"11000010100110000000000000000000"), -- -67.8 + -8.2 = -76
	(b"01000001010111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000110101100110011001100110", b"01000000111000110011001100110100"), -- 13.8 + -6.7 = 7.1
	(b"01000010011100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110000011001100110011010", b"11000010000100001100110011001110"), -- 60.6 + -96.8 = -36.2
	(b"11000010000011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011000010011001100110011", b"11000010101101111001100110011010"), -- -35.5 + -56.3 = -91.8
	(b"01000010011000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101001100000000000000000", b"11000001110101100110011001100110"), -- 56.2 + -83 = -26.8
	(b"11000010100000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101111100110011001100110", b"11000011000111111110011001100110"), -- -64.7 + -95.2 = -159.9
	(b"01000010010110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101110011001100110011", b"11000010000101001100110011001100"), -- 54.4 + -91.6 = -37.2
	(b"11000010011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110011100110011001101", b"11000011000010011011001100110011"), -- -60.8 + -76.9 = -137.7
	(b"11000001101110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000010110011001100110011", b"11000010011010000110011001100110"), -- -23.3 + -34.8 = -58.1
	(b"11000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100000000110011001100110", b"01000010011100001100110011001100"), -- -4 + 64.2 = 60.2
	(b"01000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110100100110011001100110", b"01000001111110000000000000000000"), -- 4.7 + 26.3 = 31
	(b"11000000100000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000101011001100110011010", b"11000010001001100000000000000000"), -- -4.1 + -37.4 = -41.5
	(b"11000010011001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010110100110011001100110", b"11000010111000001100110011001100"), -- -57.8 + -54.6 = -112.4
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001110101100110011001101", b"11000010001001110011001100110011"), -- 4.9 + -46.7 = -41.8
	(b"01000001101011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001010010000000000000000000", b"01000001000100011001100110011010"), -- 21.6 + -12.5 = 9.1
	(b"11000001011000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100101001100110011001101", b"01000000100100000000000000000000"), -- -14.1 + 18.6 = 4.5
	(b"01000010101000001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101011101100110011001101", b"01000011001001111011001100110100"), -- 80.3 + 87.4 = 167.7
	(b"11000010010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110000100110011001100110", b"11000001101111011001100110011010"), -- -48 + 24.3 = -23.7
	(b"01000010100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001000011001100110011010", b"01000010111011011001100110011010"), -- 78.4 + 40.4 = 118.8
	(b"11000010001111000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110011110011001100110011", b"11000010100100100000000000000000"), -- -47.1 + -25.9 = -73
	(b"11000010011011100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011000000110011001100110", b"11000000010110011001100110100000"), -- -59.5 + 56.1 = -3.4
	(b"01000010010010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000010110011001100110011", b"01000001100000000000000000000000"), -- 50.8 + -34.8 = 16
	(b"01000010100011000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001001100000000000000000", b"01000001111001011001100110011000"), -- 70.2 + -41.5 = 28.7
	(b"01000001010101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001101011011001100110011010", b"01000010000011000000000000000000"), -- 13.3 + 21.7 = 35
	(b"01000010001111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110001100110011001100110", b"01000001101110000000000000000000"), -- 47.8 + -24.8 = 23
	(b"11000000110010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010000011001100110011", b"01000010100110111001100110011001"), -- -6.3 + 84.1 = 77.8
	(b"11000001111111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000100110011001100110011", b"11000010100010001001100110011010"), -- -31.5 + -36.8 = -68.3
	(b"01000010010010000000000000000000", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"01000010010001100110011001100110"), -- 50 + -0.4 = 49.6
	(b"01000010000100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101100010110011001100110", b"01000010111110010110011001100110"), -- 36 + 88.7 = 124.7
	(b"01000010101000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100100000011001100110011", b"01000011000110001000000000000000"), -- 80.4 + 72.1 = 152.5
	(b"11000010000111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010101101100110011001101", b"01000001011000110011001100110100"), -- -39.5 + 53.7 = 14.2
	(b"01000001110101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000101001100110011001101", b"11000001001010000000000000000000"), -- 26.7 + -37.2 = -10.5
	(b"01000010000101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110011011001100110011010", b"01000010011111100000000000000000"), -- 37.8 + 25.7 = 63.5
	(b"01000010100101001100110011001101", b"00000000000000000000000000000000"),
	(b"10111110010011001100110011001101", b"01000010100101000110011001100111"), -- 74.4 + -0.2 = 74.2
	(b"01000010101000100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101001000011001100110011", b"01000011001000110011001100110011"), -- 81.1 + 82.1 = 163.2
	(b"11000010110000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101111011001100110011010", b"11000011001111110110011001100110"), -- -96.6 + -94.8 = -191.4
	(b"01000001000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101111111100110011001101", b"11000010101011100110011001100111"), -- 8.7 + -95.9 = -87.2
	(b"01000010100111101001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100111001100110011001101", b"01000010110001011100110011001101"), -- 79.3 + 19.6 = 98.9
	(b"11000010011001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010011000110011001100110", b"11000010110110001001100110011010"), -- -57.2 + -51.1 = -108.3
	(b"11000010101011110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011101010011001100110011", b"11000001110100011001100110011010"), -- -87.5 + 61.3 = -26.2
	(b"01000010100101000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001111001100110011010", b"01000011000011011110011001100110"), -- 74.1 + 67.8 = 141.9
	(b"11000010010100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101000110011001100110011", b"01000001111010001100110011001100"), -- -52.5 + 81.6 = 29.1
	(b"01000010011011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011000110011001100110011", b"01000000010000000000000000000000"), -- 59.8 + -56.8 = 3
	(b"01000010100010111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101101101100110011001101", b"01000011001000010100110011001101"), -- 69.9 + 91.4 = 161.3
	(b"11000010010001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101101011001100110011010", b"11000010100011111001100110011010"), -- -49.1 + -22.7 = -71.8
	(b"01000010101101001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101111100110011001100110", b"01000011001110011000000000000000"), -- 90.3 + 95.2 = 185.5
	(b"11000010000001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100001001001100110011010", b"11000010110001101100110011001101"), -- -33.1 + -66.3 = -99.4
	(b"11000010110000000110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"11000010101111011001100110011001"), -- -96.2 + 1.4 = -94.8
	(b"11000010101001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100010001001100110011010", b"11000011000101100100110011001101"), -- -82 + -68.3 = -150.3
	(b"11000001101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"11000001011111001100110011001101"), -- -22 + 6.2 = -15.8
	(b"01000010101100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010010000110011001100110", b"01000011000010111110011001100110"), -- 89.8 + 50.1 = 139.9
	(b"11000010000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100010110011001100110011", b"11000010110101100110011001100110"), -- -37.6 + -69.6 = -107.2
	(b"01000010101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110001100110011001100110", b"01000010100000011001100110011010"), -- 89.6 + -24.8 = 64.8
	(b"11000010100101010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100000001100110011001101", b"11000010011010011001100110011010"), -- -74.5 + 16.1 = -58.4
	(b"01000010101001100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001111100000000000000000", b"01000011000000101001100110011010"), -- 83.1 + 47.5 = 130.6
	(b"01000010010110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000000100110011001100110", b"01000001101100000000000000000000"), -- 54.6 + -32.6 = 22
	(b"01000010000111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001110101100110011001101", b"11000000111000110011001100111000"), -- 39.6 + -46.7 = -7.1
	(b"11000010000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010001001100110011010", b"11000010111101010110011001100111"), -- -38.4 + -84.3 = -122.7
	(b"01000010100100010000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110110011001100110011010", b"01000010100011011001100110011010"), -- 72.5 + -1.7 = 70.8
	(b"11000010101111010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110001010011001100110011", b"01000000011110011001100110100000"), -- -94.7 + 98.6 = 3.9
	(b"01000000100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111111100110011001101", b"11000010101101100011001100110011"), -- 4.8 + -95.9 = -91.1
	(b"11000010000011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001001111001100110011010", b"01000000110101100110011001101000"), -- -35.2 + 41.9 = 6.7
	(b"01000001010000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001011110011001100110011010", b"01000001110111011001100110011010"), -- 12.1 + 15.6 = 27.7
	(b"11000001100011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001111110100110011001100110", b"01000001010110000000000000000000"), -- -17.8 + 31.3 = 13.5
	(b"10111110010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000001100110011001100110", b"11000010000001110011001100110011"), -- -0.2 + -33.6 = -33.8
	(b"11000010001101101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110100000000000000000", b"11000010111101010110011001100110"), -- -45.7 + -77 = -122.7
	(b"11000010011000010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001001001100110011001100110", b"11000010001101111001100110011010"), -- -56.3 + 10.4 = -45.9
	(b"01000010000101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001101111001100110011001101", b"01000001010110011001100110011010"), -- 37.2 + -23.6 = 13.6
	(b"11000000101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001110100000000000000000", b"11000010010011100110011001100110"), -- -5.1 + -46.5 = -51.6
	(b"01000010101011000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001011000110011001100110", b"01000010001010111001100110011010"), -- 86 + -43.1 = 42.9
	(b"11000010101011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001010001100110011001100110", b"11000010100101100110011001100110"), -- -87.6 + 12.4 = -75.2
	(b"11000010000000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001001001100110011010", b"11000011000000100110011001100110"), -- -32.1 + -98.3 = -130.4
	(b"01000010000101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000101100110011001100110011", b"01000001111111111111111111111111"), -- 37.6 + -5.6 = 32
	(b"11000000111111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101000110011001100110", b"01000010000101001100110011001100"), -- -7.9 + 45.1 = 37.2
	(b"01000010100011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000000000110011001100110", b"01000010000111101100110011001110"), -- 71.8 + -32.1 = 39.7
	(b"01000010010100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100111101001100110011010", b"11000001110110100110011001101000"), -- 52 + -79.3 = -27.3
	(b"11000010001000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001100001000000000000000000", b"11000001101111001100110011001100"), -- -40.1 + 16.5 = -23.6
	(b"01000010101001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011001000110011001100110", b"01000001110101000000000000000000"), -- 83.6 + -57.1 = 26.5
	(b"01000010000010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001011100110011001100110011", b"01000001100111001100110011001100"), -- 34.8 + -15.2 = 19.6
	(b"11000001011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011001100000000000000000", b"11000010100100100011001100110011"), -- -15.6 + -57.5 = -73.1
	(b"01000010100100110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010110101100110011001101", b"01000011000000000110011001100110"), -- 73.7 + 54.7 = 128.4
	(b"11000010100011101001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111101100110011001100110", b"11000010110011000011001100110100"), -- -71.3 + -30.8 = -102.1
	(b"00111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101101100110011001100110", b"01000000110001100110011001100110"), -- 0.5 + 5.7 = 6.2
	(b"11000010101111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100100100011001100110011", b"11000001101100001100110011001100"), -- -95.2 + 73.1 = -22.1
	(b"01000010100101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001010001001100110011001101", b"01000010011110100000000000000001"), -- 74.8 + -12.3 = 62.5
	(b"01000010110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101111010011001100110011", b"01000011010000000011001100110011"), -- 97.6 + 94.6 = 192.2
	(b"11000010101001001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000001100110011001100110", b"11000010111001111100110011001101"), -- -82.3 + -33.6 = -115.9
	(b"11000010010111010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101111011001100110011010", b"11000001111111001100110011001100"), -- -55.3 + 23.7 = -31.6
	(b"11000010101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010011101100110011001101", b"11000010000100010011001100110011"), -- -88 + 51.7 = -36.3
	(b"11000010101011010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110111100110011001100110", b"11000010011010110011001100110011"), -- -86.6 + 27.8 = -58.8
	(b"01000010000100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000101100000000000000000", b"10111111000110011001100110000000"), -- 36.9 + -37.5 = -0.599998
	(b"11000010100110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100011110011001100110011", b"11000011000100111100110011001100"), -- -76.2 + -71.6 = -147.8
	(b"01000010100000010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111000001100110011001101", b"01000010101110010011001100110011"), -- 64.5 + 28.1 = 92.6
	(b"11000010011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"11000010011000100110011001100111"), -- -62.4 + 5.8 = -56.6
	(b"11000010101001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100010100000000000000000", b"11000001010100110011001100110000"), -- -82.2 + 69 = -13.2
	(b"11000010100111011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001001101001100110011001101", b"11000010101101000110011001100111"), -- -78.9 + -11.3 = -90.2
	(b"01000010100001001001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110111100110011001100110", b"01000010000110100000000000000001"), -- 66.3 + -27.8 = 38.5
	(b"11000010000001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100111011100110011001101", b"11000010111000000000000000000000"), -- -33.1 + -78.9 = -112
	(b"11000001101001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001001001100110011010", b"11000010101011011001100110011010"), -- -20.5 + -66.3 = -86.8
	(b"01000001001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010001100110011001100110", b"01000010011100000000000000000000"), -- 10.4 + 49.6 = 60
	(b"01000010000101010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101011110000000000000000", b"11000010010010001100110011001101"), -- 37.3 + -87.5 = -50.2
	(b"11000010000111111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010000011001100110011", b"11000010110110000000000000000000"), -- -39.9 + -68.1 = -108
	(b"11000010100100001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100000011100110011001101", b"11000011000010010011001100110100"), -- -72.3 + -64.9 = -137.2
	(b"11000010101010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101011101001100110011010", b"01000000010100110011001101000000"), -- -84 + 87.3 = 3.3
	(b"01000010100000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011001001100110011001101", b"01000001000000110011001100110100"), -- 65.4 + -57.2 = 8.2
	(b"11000010100001110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011101001100110011010", b"11000011000110101100110011001101"), -- -67.5 + -87.3 = -154.8
	(b"11000001011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101010101001100110011010", b"01000010100011010000000000000000"), -- -14.8 + 85.3 = 70.5
	(b"01000010001110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001010010110011001100110011", b"01000010000001101100110011001101"), -- 46.4 + -12.7 = 33.7
	(b"11000010001111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010001001100110011010", b"01000010000100011001100110011010"), -- -47.9 + 84.3 = 36.4
	(b"11000010100000010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101111100110011001101", b"01000001001101001100110011010000"), -- -64.6 + 75.9 = 11.3
	(b"11000001010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000000000000000000000000", b"11000001001011001100110011001101"), -- -12.8 + 2 = -10.8
	(b"01000010010000100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000111010011001100110011", b"01000010101011111001100110011010"), -- 48.5 + 39.3 = 87.8
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001010000000000000000", b"01000010011011011001100110011010"), -- -7.1 + 66.5 = 59.4
	(b"01000010101100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111100011001100110011010", b"01000010111011100110011001100110"), -- 89 + 30.2 = 119.2
	(b"01000001100010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101100011100110011001101", b"11000010100011111001100110011010"), -- 17.1 + -88.9 = -71.8
	(b"11000001000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001101101110011001100110011", b"11000010000000100000000000000000"), -- -9.6 + -22.9 = -32.5
	(b"01000001011010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010101011001100110011010", b"11000010000110101100110011001101"), -- 14.7 + -53.4 = -38.7
	(b"11000010000101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100011100011001100110011", b"01000010000001100110011001100110"), -- -37.5 + 71.1 = 33.6
	(b"11000010101001001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011111100110011001100110", b"11000001100101011001100110011100"), -- -82.3 + 63.6 = -18.7
	(b"11000010110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101100110110011001100110", b"11000011001110011011001100110011"), -- -96 + -89.7 = -185.7
	(b"11000010001101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001010000000000000000", b"11000011000100000001100110011010"), -- -45.6 + -98.5 = -144.1
	(b"01000010101101110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001101101001100110011001101", b"01000010111001001001100110011001"), -- 91.7 + 22.6 = 114.3
	(b"01000001000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101011011001100110011010", b"01000001111100011001100110011010"), -- 8.5 + 21.7 = 30.2
	(b"01000010001001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110010110011001100110011", b"01000001100000011001100110011001"), -- 41.6 + -25.4 = 16.2
	(b"01000010001111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011011010011001100110011", b"01000010110101011100110011001100"), -- 47.6 + 59.3 = 106.9
	(b"11000001101111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"11000001111000100110011001100111"), -- -23.7 + -4.6 = -28.3
	(b"11000010101110000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101001011100110011001101", b"11000011001011110000000000000000"), -- -92.1 + -82.9 = -175
	(b"01000010010011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101010011001100110011010", b"01000010001110001100110011001101"), -- 51.5 + -5.3 = 46.2
	(b"01000010101011000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101110001100110011001101", b"11000000110011001100110011010000"), -- 86 + -92.4 = -6.4
	(b"01000001100100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100011111001100110011010", b"01000010101101000011001100110100"), -- 18.3 + 71.8 = 90.1
	(b"11000001000000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101100110000000000000000", b"11000010110000110110011001100110"), -- -8.2 + -89.5 = -97.7
	(b"01000001101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001101101100110011001101", b"11000001110011011001100110011010"), -- 20 + -45.7 = -25.7
	(b"01000010101110000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011000111001100110011010", b"01000011000101010000000000000000"), -- 92.1 + 56.9 = 149
	(b"11000001100101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001010011001100110011", b"01000010001111101100110011001100"), -- -18.9 + 66.6 = 47.7
	(b"11000010010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100011010110011001100110", b"01000001101010001100110011001100"), -- -49.6 + 70.7 = 21.1
	(b"11000010101011010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100111001100110011001101", b"11000011001001010000000000000000"), -- -86.6 + -78.4 = -165
	(b"11000010100001111100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100100000000000000000000", b"11000010011111011001100110011010"), -- -67.9 + 4.5 = -63.4
	(b"01000010100010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110110000000000000000", b"01000011000100100001100110011010"), -- 68.6 + 77.5 = 146.1
	(b"01000010110001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100100110011001100110011", b"01000010101110111001100110011010"), -- 98.4 + -4.6 = 93.8
	(b"11000010101110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101000001100110011001101", b"11000010111000001001100110011001"), -- -92.2 + -20.1 = -112.3
	(b"01000010101001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101000101001100110011010", b"00111111101001100110011001000000"), -- 82.6 + -81.3 = 1.3
	(b"11000010101010100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000110010011001100110011", b"11000010001110101100110011001101"), -- -85 + 38.3 = -46.7
	(b"11000010100111111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010000000000000000000", b"11000011001000111100110011001101"), -- -79.8 + -84 = -163.8
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001100101100110011001100110", b"01000001100111011001100110011001"), -- 0.9 + 18.8 = 19.7
	(b"01000010010111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110001001100110011001101", b"01000010101000001100110011001101"), -- 55.8 + 24.6 = 80.4
	(b"01000010011011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101111001001100110011010", b"01000011000110100000000000000000"), -- 59.7 + 94.3 = 154
	(b"01000001110010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001100000110011001100110011", b"01000001000010110011001100110100"), -- 25.1 + -16.4 = 8.7
	(b"11000010100111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000000111100000000000000000000", b"11000010100011110000000000000000"), -- -79 + 7.5 = -71.5
	(b"01000010000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110000011001100110011010", b"11000010011111001100110011001110"), -- 33.6 + -96.8 = -63.2
	(b"11000010001011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101010110011001100110", b"01000010001111100110011001100110"), -- -43.1 + 90.7 = 47.6
	(b"01000010110001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011100010011001100110011", b"01000010000101111001100110011001"), -- 98.2 + -60.3 = 37.9
	(b"11000010100101010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111101100110011001100110", b"11000010110100101001100110011010"), -- -74.5 + -30.8 = -105.3
	(b"11000010100011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001010000000000000000000", b"11000010111000011001100110011010"), -- -70.8 + -42 = -112.8
	(b"01000010101011000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110001001100110011010", b"01000001000111001100110011001000"), -- 86.1 + -76.3 = 9.8
	(b"01000010001110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010011000110011001100110", b"01000010110000111001100110011010"), -- 46.7 + 51.1 = 97.8
	(b"01000010100101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001110100011001100110011010", b"01000010110010100000000000000000"), -- 74.8 + 26.2 = 101
	(b"01000010010000010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001100011001100110011010", b"01000010101110010110011001100110"), -- 48.3 + 44.4 = 92.7
	(b"01000010100110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101100011001100110011010", b"11000001010000110011001100111000"), -- 76.6 + -88.8 = -12.2
	(b"11000001100001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100111100000000000000000", b"11000010101111111100110011001101"), -- -16.9 + -79 = -95.9
	(b"01000010101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000110011001100110011010", b"01000010100101100110011001100111"), -- 84.8 + -9.6 = 75.2
	(b"11000010101100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101110100011001100110011", b"11000011001101010100110011001100"), -- -88.2 + -93.1 = -181.3
	(b"11000010001111101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110110000000000000000000", b"11000001101001011001100110011010"), -- -47.7 + 27 = -20.7
	(b"11000010001000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110001010011001100110011", b"01000010011001111001100110011001"), -- -40.7 + 98.6 = 57.9
	(b"11000000000001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100100001001100110011010", b"01000010100011000110011001100111"), -- -2.1 + 72.3 = 70.2
	(b"01000000110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011000010011001100110011", b"01000010011110101100110011001101"), -- 6.4 + 56.3 = 62.7
	(b"11000001101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111000000000000000000000", b"11000001100000011001100110011010"), -- -23.2 + 7 = -16.2
	(b"11000010100000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100000100011001100110011", b"11000011000000011100110011001100"), -- -64.7 + -65.1 = -129.8
	(b"01000000100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000011001100110011001101", b"01000001010110110011001100110100"), -- 4.9 + 8.8 = 13.7
	(b"01000010100110111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000001000000000000000000", b"01000010110111011100110011001101"), -- 77.9 + 33 = 110.9
	(b"01000001101011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110001010011001100110011", b"01000010111100001100110011001100"), -- 21.8 + 98.6 = 120.4
	(b"00111111000110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011010100110011001100110", b"01000010011011001100110011001100"), -- 0.6 + 58.6 = 59.2
	(b"01000001001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100110101001100110011010", b"01000010101011101001100110011010"), -- 10 + 77.3 = 87.3
	(b"01000010101110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001011100000000000000000000", b"01000010100110111001100110011010"), -- 92.8 + -15 = 77.8
	(b"01000001111110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101001001100110011010", b"11000010011011010011001100110100"), -- 31 + -90.3 = -59.3
	(b"01000010100110010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001001000011001100110011010", b"01000010100001001100110011001101"), -- 76.5 + -10.1 = 66.4
	(b"00000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101000110011001100110", b"11000010101101000110011001100110"), -- 0 + -90.2 = -90.2
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010100110011001100110011", b"01000010010011100110011001100110"), -- -1.2 + 52.8 = 51.6
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110010001100110011001101", b"01000001100100000000000000000000"), -- -7.1 + 25.1 = 18
	(b"11000010011011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100101111001100110011010", b"11000011000001110011001100110100"), -- -59.4 + -75.8 = -135.2
	(b"01000010000101101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010011000000000000000000", b"11000001010101001100110011001100"), -- 37.7 + -51 = -13.3
	(b"11000010011000010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010100000000000000000", b"11000011000011010100110011001101"), -- -56.3 + -85 = -141.3
	(b"11000010101101110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001100111001100110011010", b"11000010001110100110011001100110"), -- -91.5 + 44.9 = -46.6
	(b"01000010101001101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100010100110011001100110", b"01000011000110001000000000000000"), -- 83.3 + 69.2 = 152.5
	(b"00111110110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010101101100110011001101", b"11000010010101010011001100110011"), -- 0.4 + -53.7 = -53.3
	(b"01000001111101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010111001100110011001101", b"01000010101010111001100110011010"), -- 30.6 + 55.2 = 85.8
	(b"11000001011111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010010001100110011001101", b"11000010100001000011001100110011"), -- -15.9 + -50.2 = -66.1
	(b"01000010101110111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101101100000000000000000", b"01000011001110001110011001100110"), -- 93.9 + 91 = 184.9
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000111100110011001100110", b"01000010000111100000000000000000"), -- -0.1 + 39.6 = 39.5
	(b"00111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100011011100110011001101", b"11000010100010101100110011001101"), -- 1.5 + -70.9 = -69.4
	(b"01000010101100101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010001100000000000000000", b"01000010000111111001100110011010"), -- 89.4 + -49.5 = 39.9
	(b"01000010101011010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001110100110011001100110", b"01000010001000000110011001100110"), -- 86.7 + -46.6 = 40.1
	(b"11000001101010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001001101100110011001101", b"11000010011110111001100110011010"), -- -21.2 + -41.7 = -62.9
	(b"11000010011001100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001101100110011001101", b"11000010111110011100110011001101"), -- -57.5 + -67.4 = -124.9
	(b"01000010001111101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100110011001100110011010", b"01000010100001011100110011001101"), -- 47.7 + 19.2 = 66.9
	(b"11000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101110110011001100110011", b"01000010101101110011001100110011"), -- -2 + 93.6 = 91.6
	(b"01000010101010100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101101000011001100110011", b"11000000101000000000000000000000"), -- 85.1 + -90.1 = -5
	(b"11000010000100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110001100110011001100110", b"11000010011101011001100110011001"), -- -36.6 + -24.8 = -61.4
	(b"11000001110000100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100011011001100110011010", b"01000010001110100000000000000001"), -- -24.3 + 70.8 = 46.5
	(b"01000001110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001010010011001100110011", b"01000010100001010110011001100110"), -- 24.4 + 42.3 = 66.7
	(b"11000001110110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001010010110011001100110011", b"11000010000111110011001100110011"), -- -27.1 + -12.7 = -39.8
	(b"01000001100110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000010110011001100110", b"01000010111001111001100110011001"), -- 19.1 + 96.7 = 115.8
	(b"11000010101110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011011111001100110011010", b"11000011000110011000000000000000"), -- -93.6 + -59.9 = -153.5
	(b"11000010100001110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101111000000000000000000", b"01000001110100100110011001101000"), -- -67.7 + 94 = 26.3
	(b"01000001100011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111000011001100110011010", b"11000001001001100110011001101000"), -- 17.8 + -28.2 = -10.4
	(b"01000010101010000110011001100110", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"01000010101001011100110011001100"), -- 84.2 + -1.3 = 82.9
	(b"11000010100000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000000100001100110011001100110", b"11000010011101001100110011001101"), -- -65.4 + 4.2 = -61.2
	(b"01000001001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000011000110011001100110", b"01000010001110001100110011001100"), -- 11.1 + 35.1 = 46.2
	(b"11000010100011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001111000110011001100110", b"11000010111011010110011001100110"), -- -71.6 + -47.1 = -118.7
	(b"01000010010010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100101111001100110011010", b"11000001110011001100110011001110"), -- 50.2 + -75.8 = -25.6
	(b"01000010011101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000010011001100110011", b"01000000100111001100110011010000"), -- 61.2 + -56.3 = 4.9
	(b"11000001101011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011011001100110011001101", b"01000010000101100000000000000000"), -- -21.7 + 59.2 = 37.5
	(b"01000000111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100001011100110011001101", b"11000010011011100000000000000000"), -- 7.4 + -66.9 = -59.5
	(b"01000010000110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000101110011001100110011010", b"01000010001100011001100110011001"), -- 38.6 + 5.8 = 44.4
	(b"11000010100110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110100110011001100110011", b"11000010110100000000000000000000"), -- -77.6 + -26.4 = -104
	(b"01000010100001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100100000000000000000000", b"11000000101110011001100110100000"), -- 66.2 + -72 = -5.8
	(b"11000001101110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001010100011001100110011010", b"11000001000111100110011001100110"), -- -23 + 13.1 = -9.9
	(b"11000001111111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000100100000000000000000", b"01000000101000000000000000000000"), -- -31.5 + 36.5 = 5
	(b"01000010000010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100011010110011001100110", b"01000010110100100011001100110011"), -- 34.4 + 70.7 = 105.1
	(b"11000010100100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100111000000000000000000", b"11000011000101111100110011001101"), -- -73.8 + -78 = -151.8
	(b"11000010001010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100110101001100110011010", b"11000010111100000110011001100111"), -- -42.9 + -77.3 = -120.2
	(b"11000010100010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011101000000000000000000", b"11000000111011001100110011010000"), -- -68.4 + 61 = -7.4
	(b"11000010001101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001010011100110011001100110", b"11000010011010101100110011001100"), -- -45.8 + -12.9 = -58.7
	(b"01000010010110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001010000000000000000000", b"01000010110000010011001100110011"), -- 54.6 + 42 = 96.6
	(b"01000010000110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001100000011001100110011010", b"01000001101100011001100110011010"), -- 38.4 + -16.2 = 22.2
	(b"11000010100110011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010101100000000000000000", b"11000011000000100110011001100110"), -- -76.9 + -53.5 = -130.4
	(b"01000001100101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001001110011001100110011", b"11000001101110001100110011001100"), -- 18.7 + -41.8 = -23.1
	(b"01000010101011000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000011110011001100110011", b"01000010111100111100110011001100"), -- 86.1 + 35.8 = 121.9
	(b"11000001101001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000010100110011001100110011", b"11000001110000000000000000000000"), -- -20.7 + -3.3 = -24
	(b"11000010100010100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001100011001100110011010", b"11000001110001001100110011001100"), -- -69 + 44.4 = -24.6
	(b"11000001100011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000000101111001100110011001101", b"11000001001110011001100110011010"), -- -17.5 + 5.9 = -11.6
	(b"11000010101110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100000011001100110011010", b"11000011000111100110011001100110"), -- -93.6 + -64.8 = -158.4
	(b"01000010000110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000000111010011001100110011010", b"01000010001110000000000000000000"), -- 38.7 + 7.3 = 46
	(b"11000001001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100010010000000000000000", b"01000010011010000110011001100110"), -- -10.4 + 68.5 = 58.1
	(b"01000001111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001111111110011001100110011", b"10111111110000000000000000000000"), -- 30.4 + -31.9 = -1.5
	(b"01000001100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101000000000000000000000", b"11000010011101000000000000000000"), -- 19 + -80 = -61
	(b"11000010100101001001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110110001100110011001101", b"11000010110010101100110011001101"), -- -74.3 + -27.1 = -101.4
	(b"11000001000001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"11000001010010011001100110011010"), -- -8.3 + -4.3 = -12.6
	(b"01000010101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010000000000000000000000", b"01000010001001100110011001100110"), -- 89.6 + -48 = 41.6
	(b"11000001110110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001010110000000000000000000", b"11000010001000100110011001100110"), -- -27.1 + -13.5 = -40.6
	(b"11000010101001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001101001100110011010", b"11000011001101011000000000000000"), -- -82.2 + -99.3 = -181.5
	(b"01000010010101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101001100110011001101", b"01000010110001001100110011001101"), -- 53.2 + 45.2 = 98.4
	(b"01000010001110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010011001100110011001101", b"01000010110000111001100110011010"), -- 46.6 + 51.2 = 97.8
	(b"11000010100100000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010000110011001100110", b"11000011000111000100110011001100"), -- -72.1 + -84.2 = -156.3
	(b"01000010000010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001011010000000000000000000", b"01000010010000100000000000000000"), -- 34 + 14.5 = 48.5
	(b"11000010101010101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110000110000000000000000", b"01000001010000110011001100110000"), -- -85.3 + 97.5 = 12.2
	(b"01000000101101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100111011001100110011010", b"01000010101010010000000000000000"), -- 5.7 + 78.8 = 84.5
	(b"11000001111010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001010110110011001100110011", b"11000001011110110011001100110011"), -- -29.4 + 13.7 = -15.7
	(b"11000010100100011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011101001100110011010", b"01000001011001100110011001101000"), -- -72.9 + 87.3 = 14.4
	(b"01000010101100101001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001001100110011001100110", b"01000010001111101100110011001110"), -- 89.3 + -41.6 = 47.7
	(b"11000010101001100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001101000110011001100110", b"11000010000110000000000000000000"), -- -83.1 + 45.1 = -38
	(b"01000010100011010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011001010011001100110011", b"01000001010101100110011001100100"), -- 70.7 + -57.3 = 13.4
	(b"01000010101001011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100100100110011001100110", b"01000010110010100011001100110100"), -- 82.8 + 18.3 = 101.1
	(b"01000010101101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010011000000000000000000", b"01000010001000000000000000000000"), -- 91 + -51 = 40
	(b"01000010011110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010000110011001100110", b"11000001101011110011001100110010"), -- 62.3 + -84.2 = -21.9
	(b"01000001110111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010011010000110011001100110", b"01000010101010111001100110011010"), -- 27.7 + 58.1 = 85.8
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100000100110011001100110", b"01000010011010111111111111111111"), -- -6.2 + 65.2 = 59
	(b"11000010100111001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000010011001100110011", b"11000011000111101110011001100110"), -- -78.3 + -80.6 = -158.9
	(b"11000010110000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000001100000000000000000", b"11000011000000101011001100110011"), -- -97.2 + -33.5 = -130.7
	(b"11000001111010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101111001100110011001101", b"11000000101110011001100110011000"), -- -29.4 + 23.6 = -5.8
	(b"01000010101110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001100000000000000000000", b"01000010010000001100110011001100"), -- 92.2 + -44 = 48.2
	(b"11000010000101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010110000100011001100110011", b"11000011000001101110011001100110"), -- -37.8 + -97.1 = -134.9
	(b"11000010100001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011001101100110011001101", b"11000001000001111111111111111100"), -- -66.2 + 57.7 = -8.5
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101010101001100110011010", b"11000010101000101001100110011010"), -- 4 + -85.3 = -81.3
	(b"11000001110110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100010000110011001100110", b"01000010001001001100110011001100"), -- -27 + 68.2 = 41.2
	(b"01000010101011011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010100111001100110011010", b"01000011000010111100110011001101"), -- 86.9 + 52.9 = 139.8
	(b"10111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001100111000000000000000000", b"11000001101010110011001100110011"), -- -1.9 + -19.5 = -21.4
	(b"11000010010010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101000001100110011001101", b"01000001111100001100110011001110"), -- -50.3 + 80.4 = 30.1
	(b"01000010100011111001100110011010", b"00000000000000000000000000000000"),
	(b"11000001111100011001100110011010", b"01000010001001100110011001100111"), -- 71.8 + -30.2 = 41.6
	(b"11000010101000010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110000011001100110011010", b"11000010110100010110011001100110"), -- -80.5 + -24.2 = -104.7
	(b"11000010001110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011010010011001100110011", b"11000010110100010000000000000000"), -- -46.2 + -58.3 = -104.5
	(b"11000010010111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000010100000000000000000", b"11000001101001110011001100110100"), -- -55.4 + 34.5 = -20.9
	(b"11000001101110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100011011100110011001101", b"01000010001111100110011001100111"), -- -23.3 + 70.9 = 47.6
	(b"11000010100001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100010110011001100110011", b"11000010010001100110011001100110"), -- -67 + 17.4 = -49.6
	(b"11000010010000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001011100110011001100110011", b"11000010000001000000000000000000"), -- -48.2 + 15.2 = -33
	(b"11000010010111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001000011001100110011010", b"11000010110000000011001100110100"), -- -55.7 + -40.4 = -96.1
	(b"01000010001000100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101011110110011001100110", b"01000011000000000011001100110011"), -- 40.5 + 87.7 = 128.2
	(b"11000001111011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011011100000000000000000", b"11000010101100100011001100110011"), -- -29.6 + -59.5 = -89.1
	(b"11000010100001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110101011001100110011010", b"11000010101110100011001100110100"), -- -66.4 + -26.7 = -93.1
	(b"11000010101100010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101011100110011001100110", b"10111111110000000000000000000000"), -- -88.7 + 87.2 = -1.5
	(b"01000010100001010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001111101100110011001101", b"01000001100101100110011001100110"), -- 66.5 + -47.7 = 18.8
	(b"01000010000100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001111100110011001100110011", b"01000000110011001100110011001100"), -- 36.8 + -30.4 = 6.4
	(b"11000010100111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000110111001100110011010", b"11000010111010110110011001100111"), -- -78.8 + -38.9 = -117.7
	(b"11000001000111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000100111001100110011001101", b"11000000100111111111111111111111"), -- -9.9 + 4.9 = -5
	(b"01000010001101111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100110000011001100110011", b"01000010111101000000000000000000"), -- 45.9 + 76.1 = 122
	(b"01000001110010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010000101100110011001101", b"01000010100101000011001100110011"), -- 25.4 + 48.7 = 74.1
	(b"11000010000000100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100000000011001100110011", b"01000001111111001100110011001100"), -- -32.5 + 64.1 = 31.6
	(b"11000010101011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000111111001100110011010", b"11000010111111110000000000000000"), -- -87.6 + -39.9 = -127.5
	(b"01000001001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011111000110011001100110", b"01000010100100110000000000000000"), -- 10.4 + 63.1 = 73.5
	(b"01000001101110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000010000000000000000", b"11000010011001011001100110011010"), -- 23.1 + -80.5 = -57.4
	(b"11000010010001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011111100000000000000000", b"11000010111000100110011001100110"), -- -49.7 + -63.5 = -113.2
	(b"11000010001111010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010111001100110011010", b"11000011000001010001100110011010"), -- -47.3 + -85.8 = -133.1
	(b"11000010101111110110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110000011001100110011010", b"11000010100011110000000000000000"), -- -95.7 + 24.2 = -71.5
	(b"01000010101000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110110001100110011001101", b"01000010010101100110011001100110"), -- 80.7 + -27.1 = 53.6
	(b"01000010000011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110010000000000000000", b"01000010110111110011001100110011"), -- 35.1 + 76.5 = 111.6
	(b"01000010011101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101010101100110011001101", b"01000011000100110011001100110011"), -- 61.8 + 85.4 = 147.2
	(b"11000010101010011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001001101100110011001100110", b"11000010110000001001100110011010"), -- -84.9 + -11.4 = -96.3
	(b"01000001100111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100111011100110011001101", b"01000010110001010000000000000000"), -- 19.6 + 78.9 = 98.5
	(b"01000010001011010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101010000000000000000000", b"01000001101100100110011001100110"), -- 43.3 + -21 = 22.3
	(b"01000010101000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100010011001100110011010", b"01000011000101100100110011001101"), -- 81.5 + 68.8 = 150.3
	(b"01000001011010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100101011100110011001101", b"11000010011100011001100110011010"), -- 14.5 + -74.9 = -60.4
	(b"01000010101000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111010011001100110011010", b"01000010010100001100110011001101"), -- 81.4 + -29.2 = 52.2
	(b"11000001000001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100110100011001100110011", b"11000010101010110000000000000000"), -- -8.4 + -77.1 = -85.5
	(b"11000010100100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001111010100110011001100110", b"11000010110010110000000000000000"), -- -72.2 + -29.3 = -101.5
	(b"11000010101101111100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000000100000000000000000", b"11000010111110001100110011001101"), -- -91.9 + -32.5 = -124.4
	(b"11000010100110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100010011001100110011010", b"11000010011011110011001100110011"), -- -77 + 17.2 = -59.8
	(b"01000010101100000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010110110011001100110011", b"01000010000001010011001100110011"), -- 88.1 + -54.8 = 33.3
	(b"11000010100011000011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100010100000000000000000", b"11000011000010110001100110011010"), -- -70.1 + -69 = -139.1
	(b"01000010010011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101101110000000000000000", b"01000011000011101011001100110011"), -- 51.2 + 91.5 = 142.7
	(b"01000010100001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001101001001100110011001101", b"01000010001101011001100110011010"), -- 66 + -20.6 = 45.4
	(b"01000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000101100110011001100110", b"11000010000001110011001100110011"), -- 3.8 + -37.6 = -33.8
	(b"01000010001000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110001011001100110011010", b"01000010100000010110011001100110"), -- 40 + 24.7 = 64.7
	(b"01000001101010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110110011001100110011", b"01000001001110011001100110011001"), -- 21.3 + -9.7 = 11.6
	(b"11000010011110100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001101001100110011010", b"11000011000000011100110011001101"), -- -62.5 + -67.3 = -129.8
	(b"11000010100101101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100110110011001100110011", b"11000011000110010000000000000000"), -- -75.4 + -77.6 = -153
	(b"11000010001111010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010111100110011001101", b"11000011000001010011001100110011"), -- -47.3 + -85.9 = -133.2
	(b"11000010101100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101111011100110011001101", b"11000011001101110001100110011010"), -- -88.2 + -94.9 = -183.1
	(b"11000001101000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111100001100110011001101", b"11000010010010000110011001100110"), -- -20 + -30.1 = -50.1
	(b"01000001011011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011111001100110011001101", b"01000010100111000011001100110011"), -- 14.9 + 63.2 = 78.1
	(b"01000001101101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000110000110011001100110", b"11000001011100110011001100110010"), -- 22.9 + -38.1 = -15.2
	(b"11000010001011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001011111100110011001100110", b"11000001110110100110011001100111"), -- -43.2 + 15.9 = -27.3
	(b"01000010001011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011011010011001100110011", b"11000001011111001100110011001100"), -- 43.5 + -59.3 = -15.8
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101110010011001100110011", b"01000010101100100000000000000000"), -- -3.6 + 92.6 = 89
	(b"01000010101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101110100110011001100110", b"01000011001100111001100110011010"), -- 86.4 + 93.2 = 179.6
	(b"11000000011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101110011100110011001101", b"11000010110000010110011001100111"), -- -3.8 + -92.9 = -96.7
	(b"01000010011010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001001100011001100110011010", b"01000010100010101001100110011010"), -- 58.2 + 11.1 = 69.3
	(b"11000000011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010111000000000000000000", b"01000010010011011001100110011010"), -- -3.6 + 55 = 51.4
	(b"01000001011100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100101011001100110011010", b"11000000011011001100110011010000"), -- 15 + -18.7 = -3.7
	(b"01000010100001101001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000000011001100110011", b"11000001010011001100110011001000"), -- 67.3 + -80.1 = -12.8
	(b"11000010011111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100001010011001100110011", b"01000000001011001100110011000000"), -- -63.9 + 66.6 = 2.7
	(b"01000010001110000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011010110011001100110011", b"01000001111110110011001100110010"), -- 46.1 + -14.7 = 31.4
	(b"01000010001000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110110100110011001100110", b"01000001010010110011001100110100"), -- 40 + -27.3 = 12.7
	(b"11000001100001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001010000110011001100110011", b"11000000100010011001100110011010"), -- -16.5 + 12.2 = -4.3
	(b"11000010010110101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001101011110011001100110011", b"11000010100110010011001100110011"), -- -54.7 + -21.9 = -76.6
	(b"11000010011100101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101010011001100110011", b"11000001011101100110011001101000"), -- -60.7 + 45.3 = -15.4
	(b"11000010011100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001011001100110011010", b"01000001101011110011001100110100"), -- -60.9 + 82.8 = 21.9
	(b"01000000000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010100111001100110011010", b"11000010010010111001100110011010"), -- 2 + -52.9 = -50.9
	(b"01000001100110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101110001100110011001101", b"01000010110111111001100110011010"), -- 19.4 + 92.4 = 111.8
	(b"11000010100001100000000000000000", b"00000000000000000000000000000000"),
	(b"10111111101001100110011001100110", b"11000010100010001001100110011010"), -- -67 + -1.3 = -68.3
	(b"01000010000010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110111001100110011001101", b"01000010011101110011001100110100"), -- 34.2 + 27.6 = 61.8
	(b"11000010010110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011001001100110011001101", b"01000000001011001100110011010000"), -- -54.5 + 57.2 = 2.7
	(b"01000000100100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001111100110011001100110", b"01000010010100001100110011001100"), -- 4.6 + 47.6 = 52.2
	(b"11000010001000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000010010000111001100110011010"), -- -40.4 + -8.5 = -48.9
	(b"01000010101010100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010101010011001100110011", b"01000001111111100110011001100110"), -- 85.1 + -53.3 = 31.8
	(b"01000010010101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110010110011001100110", b"01000011000000100100110011001100"), -- 53.6 + 76.7 = 130.3
	(b"01000010011111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001101100110011001100110", b"01000001100100001100110011001110"), -- 63.7 + -45.6 = 18.1
	(b"11000001010101100110011001100110", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000001010111001100110011001100"), -- -13.4 + -0.4 = -13.8
	(b"11000010110001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101110100110011001100110", b"11000000110011001100110011010000"), -- -99.6 + 93.2 = -6.4
	(b"11000010100000100011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000010100100110011001100110011"), -- -65.1 + -8.5 = -73.6
	(b"01000010011100101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000100110011001100110", b"01000000100000110011001100111000"), -- 60.7 + -56.6 = 4.1
	(b"01000010100001001001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100001100110011001100110", b"01000010011110000110011001100111"), -- 66.3 + -4.2 = 62.1
	(b"01000010101111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001101001100110011001101", b"01000010010010001100110011001101"), -- 95.4 + -45.2 = 50.2
	(b"11000001110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101111111001100110011010", b"01000010100011000110011001100111"), -- -25.6 + 95.8 = 70.2
	(b"01000001110100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001101111000000000000000000", b"01000010010001101100110011001101"), -- 26.2 + 23.5 = 49.7
	(b"01000001001010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000100000000000000000000000", b"01000000110100110011001100110100"), -- 10.6 + -4 = 6.6
	(b"01000010100000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001101110001100110011001101", b"01000010001001010011001100110100"), -- 64.4 + -23.1 = 41.3
	(b"11000010100001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001001110011001100110011010", b"11000010010111000000000000000000"), -- -66.6 + 11.6 = -55
	(b"11000010010110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001100100000000000000000", b"11000001001000110011001100110100"), -- -54.7 + 44.5 = -10.2
	(b"11000001110010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011011010011001100110011", b"01000010000010000000000000000000"), -- -25.3 + 59.3 = 34
	(b"11000010000100100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000100110011001100110011", b"11000010100100101001100110011010"), -- -36.5 + -36.8 = -73.3
	(b"01000001101101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100000001001100110011010", b"11000010001001100000000000000001"), -- 22.8 + -64.3 = -41.5
	(b"11000010010101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101010010110011001100110", b"11000011000010101000000000000000"), -- -53.8 + -84.7 = -138.5
	(b"11000010000111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001010101100110011001101", b"11000010101001010000000000000000"), -- -39.8 + -42.7 = -82.5
	(b"11000010101110010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010001110011001100110011", b"11000010001010111001100110011001"), -- -92.7 + 49.8 = -42.9
	(b"01000010100010001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101001100000000000000000", b"11000001011010110011001100110000"), -- 68.3 + -83 = -14.7
	(b"11000010100101111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101101100011001100110011", b"01000001011100110011001100110000"), -- -75.9 + 91.1 = 15.2
	(b"11000010011001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100010000000000000000000", b"11000010111110110110011001100110"), -- -57.7 + -68 = -125.7
	(b"11000010010101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001000111001100110011001101", b"11000010011111100110011001100110"), -- -53.8 + -9.8 = -63.6
	(b"11000001100110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"11000001101101011001100110011001"), -- -19.3 + -3.4 = -22.7
	(b"01000001100001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000001000000000000000000", b"01000010010001100000000000000000"), -- 16.5 + 33 = 49.5
	(b"01000010101000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000001000000000000000000000", b"01000010100111100011001100110011"), -- 81.6 + -2.5 = 79.1
	(b"01000010000000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"01000010000011101100110011001101"), -- 32.4 + 3.3 = 35.7
	(b"01000010000101101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111000100110011001100110", b"01000001000101100110011001101000"), -- 37.7 + -28.3 = 9.4
	(b"11000010010011010011001100110011", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"11000010010001011001100110011001"), -- -51.3 + 1.9 = -49.4
	(b"01000010110001010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101110011001100110011010", b"01000011001111111000000000000000"), -- 98.7 + 92.8 = 191.5
	(b"01000010011000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011010000000000000000000", b"10111111101100110011001101000000"), -- 56.6 + -58 = -1.4
	(b"11000010000011010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010110101100110011001101", b"01000001100110110011001100110100"), -- -35.3 + 54.7 = 19.4
	(b"01000001111000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101001000000000000000000", b"11000010010101110011001100110011"), -- 28.2 + -82 = -53.8
	(b"11000010011101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101100100110011001100110", b"11000010101010000011001100110011"), -- -61.8 + -22.3 = -84.1
	(b"11000010000000100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110000110011001100110", b"01000010001011100110011001100110"), -- -32.6 + 76.2 = 43.6
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000001000000000000000000", b"01000010001000000000000000000000"), -- 7 + 33 = 40
	(b"11000001110101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011100000110011001100110", b"11000010101011010011001100110011"), -- -26.5 + -60.1 = -86.6
	(b"11000001100111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001010100110011001100110011", b"11000000110100110011001100110010"), -- -19.8 + 13.2 = -6.6
	(b"11000010100110010000000000000000", b"00000000000000000000000000000000"),
	(b"01000001010000000000000000000000", b"11000010100000010000000000000000"), -- -76.5 + 12 = -64.5
	(b"11000010100001101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110001000000000000000000", b"01000001111101011001100110011000"), -- -67.3 + 98 = 30.7
	(b"01000001001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010001010011001100110011", b"01000010011100100000000000000000"), -- 11.2 + 49.3 = 60.5
	(b"01000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000110000000000000000000", b"01000011000000110000000000000000"), -- 93 + 38 = 131
	(b"01000001001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100010000000000000000000", b"01000001111000001100110011001101"), -- 11.1 + 17 = 28.1
	(b"01000010000101000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100010110110011001100110", b"11000010000000100110011001100110"), -- 37.1 + -69.7 = -32.6
	(b"11000010100111010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100111101001100110011010", b"00111111001100110011001110000000"), -- -78.6 + 79.3 = 0.700005
	(b"11000001011101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100111110000000000000000", b"11000010101111011001100110011010"), -- -15.3 + -79.5 = -94.8
	(b"01000010001010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010110001101100110011001101", b"01000011000011100011001100110011"), -- 42.8 + 99.4 = 142.2
	(b"11000001100101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000000110011001100110", b"01000010011101011111111111111111"), -- -18.7 + 80.2 = 61.5
	(b"01000010101111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001010110011001100110011", b"01000010010100110011001100110011"), -- 95.6 + -42.8 = 52.8
	(b"11000010100111111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000100011001100110011010", b"11000010001011011001100110011010"), -- -79.8 + 36.4 = -43.4
	(b"10111111100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001011101001100110011001101", b"11000001100001000000000000000000"), -- -1.2 + -15.3 = -16.5
	(b"11000010010101010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001110000001100110011001101", b"11000010100110101100110011001101"), -- -53.3 + -24.1 = -77.4
	(b"01000010101000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100010000000000000000000", b"01000010110001010000000000000000"), -- 81.5 + 17 = 98.5
	(b"01000001100001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000000101011001100110011001101", b"01000001001100011001100110011010"), -- 16.5 + -5.4 = 11.1
	(b"01000010010011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000001001100110011001101", b"01000010101010100000000000000000"), -- 51.8 + 33.2 = 85
	(b"11000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001010000110011001100110", b"11000010010010111001100110011001"), -- -8.8 + -42.1 = -50.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100001001100110011001101", b"11000010100001010110011001100111"), -- -0.3 + -66.4 = -66.7
	(b"01000001110001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001001100000000000000000", b"01000010100001000011001100110011"), -- 24.6 + 41.5 = 66.1
	(b"11000010101111000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001101111001100110011010", b"11000010010000010011001100110010"), -- -94.2 + 45.9 = -48.3
	(b"01000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100101100110011001101", b"11000010100001101001100110011010"), -- 6.1 + -73.4 = -67.3
	(b"11000001100011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000110111001100110011001101", b"11000001110001011001100110011001"), -- -17.8 + -6.9 = -24.7
	(b"01000010001100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010000101100110011001101", b"01000010101110101001100110011010"), -- 44.6 + 48.7 = 93.3
	(b"01000010010010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010110000001001100110011010", b"01000011000100100100110011001101"), -- 50 + 96.3 = 146.3
	(b"11000010101110110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101100110011001100110", b"11000011001110001110011001100110"), -- -93.7 + -91.2 = -184.9
	(b"11000010010101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000000000000000000000", b"11000011000001010110011001100110"), -- -53.4 + -80 = -133.4
	(b"01000010001101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000101011001100110011010", b"01000010101001100000000000000000"), -- 45.6 + 37.4 = 83
	(b"11000001001010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101110100110011001100110", b"01000001010011001100110011001100"), -- -10.5 + 23.3 = 12.8
	(b"11000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100101010000000000000000", b"11000010101001100011001100110011"), -- -8.6 + -74.5 = -83.1
	(b"01000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001111101000000000000000000", b"11000001110001110011001100110011"), -- 5.6 + -30.5 = -24.9
	(b"11000001101001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000100111001100110011001101", b"11000001110011011001100110011001"), -- -20.8 + -4.9 = -25.7
	(b"11000010011011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001010010011001100110011", b"11000001100010110011001100110100"), -- -59.7 + 42.3 = -17.4
	(b"11000001111110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001111100110011001101", b"01000010000100110011001100110100"), -- -31.1 + 67.9 = 36.8
	(b"01000010110000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001111101100110011001100110", b"01000011000000001001100110011010"), -- 97.8 + 30.8 = 128.6
	(b"01000001011101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010110000000000000000000", b"11000010000110100110011001100110"), -- 15.4 + -54 = -38.6
	(b"11000010000100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000011111001100110011010", b"11000010100100011001100110011010"), -- -36.9 + -35.9 = -72.8
	(b"01000001100000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001101100110011001100110", b"01000010011101110011001100110011"), -- 16.2 + 45.6 = 61.8
	(b"01000001011010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011000000000000000000000", b"01000010100011010110011001100110"), -- 14.7 + 56 = 70.7
	(b"01000010001101001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000011000000000000000000", b"01000001001000110011001100110100"), -- 45.2 + -35 = 10.2
	(b"11000010000111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100000000000000000000", b"11000010000001010011001100110011"), -- -39.8 + 6.5 = -33.3
	(b"11000010100000000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010000101100110011001101", b"11000001011101100110011001100100"), -- -64.1 + 48.7 = -15.4
	(b"01000010000000100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011110011001100110011", b"11000010010111000110011001100110"), -- 32.5 + -87.6 = -55.1
	(b"01000010100011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000101001100110011001101", b"01000010110110001100110011001100"), -- 71.2 + 37.2 = 108.4
	(b"11000010101110100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011010000000000000000000", b"11000010110101110110011001100110"), -- -93.2 + -14.5 = -107.7
	(b"11000010100000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101111111100110011001101", b"01000001111111011001100110011100"), -- -64.2 + 95.9 = 31.7
	(b"01000001111010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000101100000000000000000", b"11000001000001100110011001100110"), -- 29.1 + -37.5 = -8.4
	(b"11000010110001000011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110001001100110011001101", b"11000010100100110000000000000000"), -- -98.1 + 24.6 = -73.5
	(b"00111111111100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001110110011001100110", b"01000010100010110011001100110011"), -- 1.9 + 67.7 = 69.6
	(b"01000010101100101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001101000000000000000000", b"01000011000001100100110011001101"), -- 89.3 + 45 = 134.3
	(b"11000010001001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010111110011001100110011", b"11000010110000110000000000000000"), -- -41.7 + -55.8 = -97.5
	(b"01000001110001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"01000001011110000000000000000000"), -- 24.6 + -9.1 = 15.5
	(b"11000010100000100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010111101100110011001101", b"11000010111100011001100110011010"), -- -65.1 + -55.7 = -120.8
	(b"11000001010100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111111001100110011001101", b"11000010001100100110011001100110"), -- -13 + -31.6 = -44.6
	(b"11000010011010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010000010000110011001100110", b"11000010101110100000000000000000"), -- -58.9 + -34.1 = -93
	(b"11000001100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101011110011001100110011", b"11000010110101001100110011001100"), -- -18.8 + -87.6 = -106.4
	(b"01000010010010101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001100011001100110011001101", b"01000010000001000110011001100110"), -- 50.7 + -17.6 = 33.1
	(b"11000010101011011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010111000110011001100110", b"11000011000011100000000000000000"), -- -86.9 + -55.1 = -142
	(b"01000001001001100110011001100110", b"00000000000000000000000000000000"),
	(b"00111111101100110011001100110011", b"01000001001111001100110011001100"), -- 10.4 + 1.4 = 11.8
	(b"01000010101101011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001111001100110011010", b"01000011000111101011001100110100"), -- 90.9 + 67.8 = 158.7
	(b"01000001101000100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001100001100110011001101", b"01000010100000010000000000000000"), -- 20.3 + 44.2 = 64.5
	(b"11000010011000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100111101100110011001101", b"11000011000010000001100110011010"), -- -56.7 + -79.4 = -136.1
	(b"11000010010110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001011000000000000000000000", b"11000010001000100110011001100110"), -- -54.6 + 14 = -40.6
	(b"11000001000011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101000100000000000000000", b"01000010100100000011001100110011"), -- -8.9 + 81 = 72.1
	(b"01000010101011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111111100110011001100110011", b"01000010101100001001100110011010"), -- 86.4 + 1.9 = 88.3
	(b"11000010010111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010110001000110011001100110", b"01000010001011001100110011001100"), -- -55 + 98.2 = 43.2
	(b"01000010101100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001110110011001100110", b"01000011001011011000000000000000"), -- 89.8 + 83.7 = 173.5
	(b"01000010011101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111101100110011001101", b"11000010000010000000000000000000"), -- 61.4 + -95.4 = -34
	(b"10111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100110000000000000000000", b"01000010100101111100110011001101"), -- -0.1 + 76 = 75.9
	(b"01000001011000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001100010011001100110011", b"01000010011010010011001100110011"), -- 14 + 44.3 = 58.3
	(b"11000001001110110011001100110011", b"00000000000000000000000000000000"),
	(b"10111111101100110011001100110011", b"11000001010100011001100110011001"), -- -11.7 + -1.4 = -13.1
	(b"11000010001111101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111111110011001100110011", b"11000001011111001100110011001110"), -- -47.7 + 31.9 = -15.8
	(b"11000010000101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100001001001100110011010", b"11000010110100000011001100110100"), -- -37.8 + -66.3 = -104.1
	(b"01000001011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100110010110011001100110", b"11000010011101000110011001100110"), -- 15.6 + -76.7 = -61.1
	(b"01000010100111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011110110011001100110011", b"01000001011110011001100110011100"), -- 78.4 + -62.8 = 15.6
	(b"01000010100100101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000110110011001100110011", b"01000010000010100110011001100111"), -- 73.4 + -38.8 = 34.6
	(b"01000010011001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001001100110011001100110", b"01000010110001101001100110011010"), -- 57.7 + 41.6 = 99.3
	(b"11000001100010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110100011001100110011", b"01000010011011101100110011001100"), -- -17.4 + 77.1 = 59.7
	(b"01000010100010111001100110011010", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"01000010100011100011001100110100"), -- 69.8 + 1.3 = 71.1
	(b"11000010101100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000011100000000000000000", b"11000010111101111100110011001101"), -- -88.4 + -35.5 = -123.9
	(b"01000010101010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000101001100110011001101", b"01000010111100100110011001100110"), -- 84 + 37.2 = 121.2
	(b"01000010001010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001011101100110011001100110", b"01000001110101001100110011001101"), -- 42 + -15.4 = 26.6
	(b"11000001101110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000000100110011001100110011", b"11000001101001110011001100110100"), -- -23.2 + 2.3 = -20.9
	(b"10111111110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111000000000000000000", b"01000010010101100000000000000000"), -- -1.5 + 55 = 53.5
	(b"01000000110100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000110101100110011001101", b"11000010000000000110011001100111"), -- 6.6 + -38.7 = -32.1
	(b"01000010101111110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010000101100110011001101", b"01000010001110111111111111111111"), -- 95.7 + -48.7 = 47
	(b"11000010011100010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000001100000000000000000", b"11000010101110111001100110011010"), -- -60.3 + -33.5 = -93.8
	(b"01000010010110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001011100011001100110011010", b"01000010100010110000000000000000"), -- 54.4 + 15.1 = 69.5
	(b"11000010001110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100001010110011001100110", b"11000010111000110011001100110011"), -- -46.9 + -66.7 = -113.6
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010000110011001100110011", b"01000010010100110011001100110011"), -- 4 + 48.8 = 52.8
	(b"01000001101101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011100101100110011001101", b"11000010000110001100110011001101"), -- 22.5 + -60.7 = -38.2
	(b"01000010000001000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101011100110011001100110", b"01000001001101001100110011001100"), -- 33.1 + -21.8 = 11.3
	(b"11000010101000010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000010110011001100110", b"11000011001100010011001100110011"), -- -80.5 + -96.7 = -177.2
	(b"11000010110000101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100010000011001100110011", b"11000011001001011000000000000000"), -- -97.4 + -68.1 = -165.5
	(b"11000010101110111100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100110001100110011001101", b"11000010100101011001100110011010"), -- -93.9 + 19.1 = -74.8
	(b"01000001101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101110001100110011001101", b"01000010111000110011001100110100"), -- 21.2 + 92.4 = 113.6
	(b"11000010010100010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100010000011001100110011", b"01000001011111001100110011001100"), -- -52.3 + 68.1 = 15.8
	(b"11000010001101010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101000000000000000000000", b"01000010000010101100110011001101"), -- -45.3 + 80 = 34.7
	(b"11000000011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001101100110011001101", b"11000010100011011100110011001101"), -- -3.5 + -67.4 = -70.9
	(b"11000010110000000011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110001110011001100110011", b"11000010100011100110011001100110"), -- -96.1 + 24.9 = -71.2
	(b"11000010101001110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100111011100110011001101", b"11000011001000100110011001100110"), -- -83.5 + -78.9 = -162.4
	(b"01000001000101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010000111001100110011001101", b"01000010010000100110011001100110"), -- 9.4 + 39.2 = 48.6
	(b"11000010100111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011100000000000000000000", b"11000001100110011001100110011000"), -- -79.2 + 60 = -19.2
	(b"11000010011010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101101010110011001100110", b"01000010000000010011001100110010"), -- -58.4 + 90.7 = 32.3
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001010010110011001100110011", b"11000000110100000000000000000000"), -- 6.2 + -12.7 = -6.5
	(b"11000010010001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101000110011001100110", b"01000010001000100110011001100110"), -- -49.6 + 90.2 = 40.6
	(b"11000010010001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100100110110011001100110", b"01000001110001011001100110011000"), -- -49 + 73.7 = 24.7
	(b"11000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001101000000000000000000", b"11000010010011001100110011001101"), -- -6.2 + -45 = -51.2
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100011011001100110011010", b"01000010100100110011001100110100"), -- 2.8 + 70.8 = 73.6
	(b"01000010000111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100011100000000000000000", b"01000010110111010000000000000000"), -- 39.5 + 71 = 110.5
	(b"11000010100000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100111010011001100110011", b"11000011000011110100110011001100"), -- -64.7 + -78.6 = -143.3
	(b"01000001100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001100000000000000000000", b"11000001110010011001100110011010"), -- 18.8 + -44 = -25.2
	(b"11000001110100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000101100110011001101", b"11000010101001011001100110011010"), -- -26.1 + -56.7 = -82.8
	(b"01000001110101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001000110011001100110011", b"01000010100001110011001100110011"), -- 26.8 + 40.8 = 67.6
	(b"01000010011010100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001100001100110011001101", b"01000001011001001100110011001100"), -- 58.5 + -44.2 = 14.3
	(b"11000010101010111100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100000110011001100110011", b"11000010100010110000000000000000"), -- -85.9 + 16.4 = -69.5
	(b"01000010001111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100011000000000000000000", b"01000001111011000000000000000000"), -- 47 + -17.5 = 29.5
	(b"01000001101000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100110110110011001100110", b"11000010011001011111111111111111"), -- 20.2 + -77.7 = -57.5
	(b"01000010010011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010010011100000000000000000", b"01000010110011101001100110011010"), -- 51.8 + 51.5 = 103.3
	(b"01000010010000100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100011110011001100110011", b"11000001101110001100110011001100"), -- 48.5 + -71.6 = -23.1
	(b"01000001111000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101111110000000000000000", b"11000010100001101100110011001101"), -- 28.1 + -95.5 = -67.4
	(b"11000010010000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100001010000000000000000", b"11000010111001100011001100110011"), -- -48.6 + -66.5 = -115.1
	(b"11000001000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001110000000000000000000", b"11000010010110110011001100110011"), -- -8.8 + -46 = -54.8
	(b"01000010110001110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100100110110011001100110", b"01000011001011010110011001100110"), -- 99.7 + 73.7 = 173.4
	(b"01000010010011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011010000110011001100110", b"01000010110110100011001100110011"), -- 51 + 58.1 = 109.1
	(b"01000001100001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110100001100110011001101", b"11000001000110000000000000000000"), -- 16.6 + -26.1 = -9.5
	(b"01000000010000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010111011001100110011010", b"01000010011010011001100110011010"), -- 3 + 55.4 = 58.4
	(b"01000010101101100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011010110011001100110011", b"01000011000101011110011001100110"), -- 91.1 + 58.8 = 149.9
	(b"01000001111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010001011001100110011010", b"01000010101000010011001100110100"), -- 31.2 + 49.4 = 80.6
	(b"01000010110000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101110110011001100110011", b"01000011001111110001100110011010"), -- 97.5 + 93.6 = 191.1
	(b"01000001110111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010110000011001100110011010", b"11000010100010011100110011001101"), -- 27.9 + -96.8 = -68.9
	(b"11000000111000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110010011001100110011", b"01000010100010110000000000000000"), -- -7.1 + 76.6 = 69.5
	(b"11000010000101110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101111000110011001100110", b"11000011000001000000000000000000"), -- -37.8 + -94.2 = -132
	(b"11000010101001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111001011001100110011010", b"11000010010101111001100110011001"), -- -82.6 + 28.7 = -53.9
	(b"11000010010110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000101000110011001100110", b"11000010101101101100110011001100"), -- -54.3 + -37.1 = -91.4
	(b"01000001101111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001110011011001100110011010", b"01000010010001100110011001100110"), -- 23.9 + 25.7 = 49.6
	(b"01000001111101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010111101100110011001101", b"11000001110010000000000000000000"), -- 30.7 + -55.7 = -25
	(b"01000010101100010110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110011001100110011001101", b"01000010111001001001100110011001"), -- 88.7 + 25.6 = 114.3
	(b"11000010110001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101101000011001100110011", b"11000001000011100110011001101000"), -- -99 + 90.1 = -8.9
	(b"01000010010001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101001110011001100110011", b"01000011000001001100110011001101"), -- 49.2 + 83.6 = 132.8
	(b"01000001110101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100100001001100110011010", b"11000010001101100110011001100111"), -- 26.7 + -72.3 = -45.6
	(b"11000010100110100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010011100110011001100110", b"11000011000000001001100110011010"), -- -77 + -51.6 = -128.6
	(b"11000010101101100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000011001100110011001101", b"11000010111111001001100110011010"), -- -91.1 + -35.2 = -126.3
	(b"01000010001000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110001110011001100110011", b"01000011000011000100110011001101"), -- 40.7 + 99.6 = 140.3
	(b"11000010110001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000000000000000000000", b"11000011000110100110011001100110"), -- -98.4 + -56 = -154.4
	(b"11000010101101110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001010011100110011001100110", b"11000010110100010011001100110011"), -- -91.7 + -12.9 = -104.6
	(b"01000010001101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101110000000000000000000", b"01000011000010011100110011001101"), -- 45.8 + 92 = 137.8
	(b"11000010001011101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000010011001100110011010", b"11000001000101001100110011001100"), -- -43.7 + 34.4 = -9.3
	(b"11000001101010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"11000001100110000000000000000000"), -- -21.1 + 2.1 = -19
	(b"01000010011110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100100001001100110011010", b"01000011000001101011001100110100"), -- 62.4 + 72.3 = 134.7
	(b"01000001111111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010101001100110011001101", b"01000010101010010110011001100110"), -- 31.5 + 53.2 = 84.7
	(b"11000001100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100001001100110011001101", b"11000010101001100110011001100110"), -- -16.8 + -66.4 = -83.2
	(b"11000010011101111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001111001100110011001101", b"11000001011010110011001100110100"), -- -61.9 + 47.2 = -14.7
	(b"01000010110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101110101001100110011010", b"01000000001011001100110011000000"), -- 96 + -93.3 = 2.7
	(b"01000010000001010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001111001100110011001101", b"11000001010111100110011001101000"), -- 33.3 + -47.2 = -13.9
	(b"01000010101000100011001100110011", b"00000000000000000000000000000000"),
	(b"01000001010101001100110011001101", b"01000010101111001100110011001101"), -- 81.1 + 13.3 = 94.4
	(b"11000001110101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110111000000000000000000", b"11000010010110001100110011001101"), -- -26.7 + -27.5 = -54.2
	(b"01000001011100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100000010110011001100110", b"01000010100111110110011001100110"), -- 15 + 64.7 = 79.7
	(b"01000010100001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001110101001100110011001101", b"01000010101111001100110011001101"), -- 67.8 + 26.6 = 94.4
	(b"01000010001010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101101010110011001100110", b"11000010010000011111111111111111"), -- 42.2 + -90.7 = -48.5
	(b"11000010000111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100011100110011001100110", b"01000001111111011001100110011000"), -- -39.5 + 71.2 = 31.7
	(b"01000010101110000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010001000110011001100110", b"01000011000011010100110011001100"), -- 92.2 + 49.1 = 141.3
	(b"11000010100000110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101100000011001100110011", b"01000001101100110011001100110100"), -- -65.7 + 88.1 = 22.4
	(b"01000010010010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101110011001100110011", b"11000010001001000000000000000000"), -- 50.6 + -91.6 = -41
	(b"11000010101100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110100110011001100110011", b"11000010101001100000000000000000"), -- -89.6 + 6.6 = -83
	(b"11000010100001100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101110011100110011001101", b"01000001110011100110011001101000"), -- -67.1 + 92.9 = 25.8
	(b"01000000100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000111001100110011010", b"11000010101110111001100110011010"), -- 4 + -97.8 = -93.8
	(b"11000010100111101001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011101101100110011001101", b"11000011000011010000000000000000"), -- -79.3 + -61.7 = -141
	(b"01000010011011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101110101001100110011010", b"01000011000110001011001100110100"), -- 59.4 + 93.3 = 152.7
	(b"01000010100000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001000011100110011001100110", b"01000010100100100011001100110011"), -- 64.2 + 8.9 = 73.1
	(b"01000010011000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011110100000000000000000", b"11000000110011001100110011010000"), -- 56.1 + -62.5 = -6.4
	(b"01000010100011011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000110000000000000000", b"01000011001010000110011001100110"), -- 70.9 + 97.5 = 168.4
	(b"11000010101000101001100110011010", b"00000000000000000000000000000000"),
	(b"01000001010001001100110011001101", b"11000010100010100000000000000000"), -- -81.3 + 12.3 = -69
	(b"11000010010000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100101001001100110011010", b"11000010111101100011001100110100"), -- -48.8 + -74.3 = -123.1
	(b"01000010100100000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011011000110011001100110", b"01000011000000110100110011001100"), -- 72.2 + 59.1 = 131.3
	(b"01000001111001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110011100110011001101", b"01000010110100111001100110011010"), -- 28.9 + 76.9 = 105.8
	(b"01000001100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001001010110011001100110011", b"01000000110100000000000000000010"), -- 17.2 + -10.7 = 6.5
	(b"01000010110000100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000110011001100110011010", b"01000011000001111000000000000000"), -- 97.1 + 38.4 = 135.5
	(b"00111111011001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110001000000000000000000", b"01000001110010110011001100110011"), -- 0.9 + 24.5 = 25.4
	(b"11000010001010111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100111000000000000000000", b"11000001101110110011001100110100"), -- -42.9 + 19.5 = -23.4
	(b"11000010101100100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100011000110011001100110", b"11000011000111110100110011001100"), -- -89.1 + -70.2 = -159.3
	(b"11000010100011010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000010000000000000000000", b"11000010100111100110011001100110"), -- -70.7 + -8.5 = -79.2
	(b"01000010011110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101110010011001100110011", b"11000001111100011001100110011000"), -- 62.4 + -92.6 = -30.2
	(b"11000010100010110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000000111001100110011010", b"11000010110011001100110011001101"), -- -69.5 + -32.9 = -102.4
	(b"01000010100101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110111110011001100110011", b"01000010001110111001100110011010"), -- 74.8 + -27.9 = 46.9
	(b"11000010101000110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110001100000000000000000", b"01000001100010100110011001101000"), -- -81.7 + 99 = 17.3
	(b"11000010011110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101101110011001100110011", b"01000001111010110011001100110010"), -- -62.2 + 91.6 = 29.4
	(b"01000001101111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000000011001100110011", b"01000010110011111001100110011010"), -- 23.7 + 80.1 = 103.8
	(b"11000010101110100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101000010000000000000000", b"11000001010010000000000000000000"), -- -93 + 80.5 = -12.5
	(b"01000001011001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100011001001100110011010", b"01000010101010010011001100110100"), -- 14.3 + 70.3 = 84.6
	(b"11000001111111110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101110011001100110011010", b"11000010000101101100110011001101"), -- -31.9 + -5.8 = -37.7
	(b"01000010110000100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010010000110011001100110", b"01000011000100110100110011001100"), -- 97.2 + 50.1 = 147.3
	(b"11000001001000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000001001100110011001100110", b"11000000111100110011001100110011"), -- -10.2 + 2.6 = -7.6
	(b"01000010100000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101100011001100110011", b"11000001110100110011001100110100"), -- 64.7 + -91.1 = -26.4
	(b"11000001101001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000100000000000000000000", b"01000001011101100110011001100110"), -- -20.6 + 36 = 15.4
	(b"01000010001100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001001111100110011001100110", b"01000010011000000110011001100110"), -- 44.2 + 11.9 = 56.1
	(b"01000001101001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110010011001100110011010", b"01000001011001100110011001100111"), -- 20.7 + -6.3 = 14.4
	(b"01000010100100111100110011001101", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"01000010100001000011001100110011"), -- 73.9 + -7.8 = 66.1
	(b"11000010100100010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100011101100110011001101", b"11000011000011111110011001100110"), -- -72.5 + -71.4 = -143.9
	(b"11000010100101011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101011010110011001100110", b"01000001001111001100110011001000"), -- -74.9 + 86.7 = 11.8
	(b"11000000100011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101010111001100110011010", b"11000010101101000110011001100111"), -- -4.4 + -85.8 = -90.2
	(b"01000010100100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011110010011001100110011", b"01000001001000011001100110011100"), -- 72.4 + -62.3 = 10.1
	(b"01000010000110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100001001100110011001101", b"01000010110100010011001100110100"), -- 38.2 + 66.4 = 104.6
	(b"01000010101111001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010110001011100110011001101", b"01000011010000010011001100110100"), -- 94.3 + 98.9 = 193.2
	(b"11000010100110000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101000000011001100110011", b"01000000100000000000000000000000"), -- -76.1 + 80.1 = 4
	(b"01000010101001110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101110000000000000000000", b"11000001000001001100110011010000"), -- 83.7 + -92 = -8.3
	(b"01000001010111001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"01000001011110000000000000000000"), -- 13.8 + 1.7 = 15.5
	(b"01000010101010000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101000000000000000000", b"01000011000111100001100110011010"), -- 84.1 + 74 = 158.1
	(b"01000010101111101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101110101001100110011010", b"01000011001111001001100110011010"), -- 95.3 + 93.3 = 188.6
	(b"00111101110011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101111101100110011001101", b"11000010101111101001100110011010"), -- 0.1 + -95.4 = -95.3
	(b"11000010000010101100110011001101", b"00000000000000000000000000000000"),
	(b"10111110110011001100110011001101", b"11000010000011000110011001100111"), -- -34.7 + -0.4 = -35.1
	(b"01000000110001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101000110011001100110011", b"01000010101011111001100110011001"), -- 6.2 + 81.6 = 87.8
	(b"11000010001100000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010011001010011001100110011", b"11000010110010101100110011001100"), -- -44.1 + -57.3 = -101.4
	(b"01000010101000011100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110110011001100110011010", b"01000010010101101100110011001101"), -- 80.9 + -27.2 = 53.7
	(b"11000010101101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010101010110011001100110011", b"11000000110000000000000000000000"), -- -91.6 + 85.6 = -6
	(b"01000010000000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001100000000000000000000", b"01000010100110000011001100110011"), -- 32.1 + 44 = 76.1
	(b"01000001110111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010110000110000000000000000", b"01000010111110101100110011001101"), -- 27.9 + 97.5 = 125.4
	(b"11000010001101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100001111100110011001101", b"11000010111000011100110011001101"), -- -45 + -67.9 = -112.9
	(b"01000010101110001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000010110011001100110011010", b"01000010101100100000000000000000"), -- 92.4 + -3.4 = 89
	(b"11000010101101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110001110000000000000000", b"01000001000100011001100110011000"), -- -90.4 + 99.5 = 9.1
	(b"11000010000010101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100111011100110011001101", b"11000010111000110011001100110100"), -- -34.7 + -78.9 = -113.6
	(b"11000010010101111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101101000110011001100110", b"11000011000100000001100110011010"), -- -53.9 + -90.2 = -144.1
	(b"01000010100010100011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010011011001100110011010", b"01000001100011011001100110011000"), -- 69.1 + -51.4 = 17.7
	(b"01000010100101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100101110011001100110011", b"01000010101110111100110011001101"), -- 75 + 18.9 = 93.9
	(b"11000001011011001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111101001100110011001100110", b"11000001010110000000000000000000"), -- -14.8 + 1.3 = -13.5
	(b"01000010011100000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011100011001100110011010", b"01000010111100010000000000000000"), -- 60.1 + 60.4 = 120.5
	(b"01000001101100001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011101010011001100110011", b"11000010000111001100110011001100"), -- 22.1 + -61.3 = -39.2
	(b"11000010001000111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100100000000000000000000", b"11000001101101110011001100110100"), -- -40.9 + 18 = -22.9
	(b"11000010011010101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010011000110011001100110011", b"10111111111100110011001101000000"), -- -58.7 + 56.8 = -1.9
	(b"01000001111011011001100110011010", b"00000000000000000000000000000000"),
	(b"01000000111000110011001100110011", b"01000010000100110011001100110011"), -- 29.7 + 7.1 = 36.8
	(b"01000010110001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100001101001100110011010", b"01000010000000000110011001100110"), -- 99.4 + -67.3 = 32.1
	(b"11000010101000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100010101100110011001101", b"11000001001100000000000000000000"), -- -80.4 + 69.4 = -11
	(b"11000010001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100111110000000000000000", b"01000010000010101100110011001101"), -- -44.8 + 79.5 = 34.7
	(b"01000010100101010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010001011001100110011010", b"01000010111101111100110011001101"), -- 74.5 + 49.4 = 123.9
	(b"01000010100001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001110000100110011001100110", b"01000010101101001001100110011010"), -- 66 + 24.3 = 90.3
	(b"01000010110000100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110100100110011001100110", b"01000010111101110000000000000000"), -- 97.2 + 26.3 = 123.5
	(b"01000001111111000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001010110011001100110011", b"11000001001101001100110011001100"), -- 31.5 + -42.8 = -11.3
	(b"11000010010010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001100010000000000000000000", b"11000010100001100000000000000000"), -- -50 + -17 = -67
	(b"01000010101110000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010110001000011001100110011", b"01000011001111100001100110011010"), -- 92 + 98.1 = 190.1
	(b"11000010001100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100010111001100110011010", b"11000010111001010011001100110100"), -- -44.8 + -69.8 = -114.6
	(b"01000010011110010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001010100000000000000000", b"01000010110100011001100110011010"), -- 62.3 + 42.5 = 104.8
	(b"11000010101011010000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101101001100110011001101", b"01000000011110011001100110100000"), -- -86.5 + 90.4 = 3.9
	(b"01000010101001101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001100101000000000000000000", b"01000010100000011100110011001101"), -- 83.4 + -18.5 = 64.9
	(b"11000010100110100011001100110011", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000010100110010000000000000000"), -- -77.1 + 0.6 = -76.5
	(b"11000001100100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101000000000000000000", b"11000010110110001001100110011010"), -- -18.3 + -90 = -108.3
	(b"01000001101111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111111100110011001101", b"11000010100100000110011001100110"), -- 23.7 + -95.9 = -72.2
	(b"01000010000011101100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001110110011001100110011", b"11000001001100011001100110011000"), -- 35.7 + -46.8 = -11.1
	(b"01000010000100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001011111001100110011001101", b"01000010010100100110011001100110"), -- 36.8 + 15.8 = 52.6
	(b"01000010010011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010000010011001100110011", b"01000000010001100110011001110000"), -- 51.4 + -48.3 = 3.1
	(b"01000010000101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010101001100110011001101", b"01000010101101010011001100110100"), -- 37.4 + 53.2 = 90.6
	(b"11000010000101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000000000001100110011001100110", b"11000010000011000110011001100111"), -- -37.2 + 2.1 = -35.1
	(b"11000010001101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101100001100110011001101", b"01000010001011001100110011001101"), -- -45.2 + 88.4 = 43.2
	(b"11000010011011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001001111001100110011010", b"11000001100010011001100110011000"), -- -59.1 + 41.9 = -17.2
	(b"11000001100001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101000010110011001100110", b"01000010100000000011001100110011"), -- -16.6 + 80.7 = 64.1
	(b"01000010100101100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101100101001100110011010", b"01000011001001000100110011001101"), -- 75 + 89.3 = 164.3
	(b"11000001100111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001001001001100110011001101", b"11000001111100000000000000000000"), -- -19.7 + -10.3 = -30
	(b"11000001110110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101110000000000000000", b"11000010111011010000000000000000"), -- -27 + -91.5 = -118.5
	(b"01000010010010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110000011001100110011010", b"01000001110100011001100110011010"), -- 50.4 + -24.2 = 26.2
	(b"01000010110000011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010100111110011001100110011", b"01000001100010100110011001101000"), -- 96.9 + -79.6 = 17.3
	(b"01000001100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001011100110011001100110011", b"00111111010011001100110011010000"), -- 16 + -15.2 = 0.8
	(b"11000001100000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100100001100110011001101", b"01000010011000010011001100110100"), -- -16.1 + 72.4 = 56.3
	(b"01000010100100011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000011001100110011010", b"11000000111111001100110011010000"), -- 72.9 + -80.8 = -7.9
	(b"01000010100001010110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111011001100110011001101", b"01000010011011010011001100110010"), -- 66.7 + -7.4 = 59.3
	(b"01000010000110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100000100110011001100110", b"01000010010111000000000000000000"), -- 38.7 + 16.3 = 55
	(b"11000010100000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011010000000000000000000", b"11000010100111010110011001100110"), -- -64.2 + -14.5 = -78.7
	(b"01000010010000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101001001100110011001101", b"01000010100010101100110011001101"), -- 48.8 + 20.6 = 69.4
	(b"01000010101010100110011001100110", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"01000010100110110011001100110011"), -- 85.2 + -7.6 = 77.6
	(b"11000010100010001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001111111001100110011010", b"11000001101000110011001100110100"), -- -68.3 + 47.9 = -20.4
	(b"11000010100010010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000011100110011001100110", b"11000010110100000011001100110011"), -- -68.5 + -35.6 = -104.1
	(b"01000000101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100110100000000000000000", b"01000010101001000110011001100110"), -- 5.2 + 77 = 82.2
	(b"01000010010111100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011100000000000000000000", b"01000010001000100110011001100110"), -- 55.6 + -15 = 40.6
	(b"01000010101011011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000101001100110011001101", b"01000010010001101100110011001101"), -- 86.9 + -37.2 = 49.7
	(b"11000010101000000110011001100110", b"00000000000000000000000000000000"),
	(b"00111111011001100110011001100110", b"11000010100111101001100110011001"), -- -80.2 + 0.9 = -79.3
	(b"11000010011010100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011110100110011001100110", b"01000000100000000000000000000000"), -- -58.6 + 62.6 = 4
	(b"01000010101100010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101101000011001100110011", b"01000011001100101100110011001100"), -- 88.7 + 90.1 = 178.8
	(b"11000010100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001111010011001100110011", b"11000010110111101001100110011010"), -- -64 + -47.3 = -111.3
	(b"10111111100000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101101000011001100110011", b"11000010101101100011001100110011"), -- -1 + -90.1 = -91.1
	(b"01000001111110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001000111100110011001100110", b"01000010001001000110011001100110"), -- 31.2 + 9.9 = 41.1
	(b"01000010110001101100110011001101", b"00000000000000000000000000000000"),
	(b"01000000110001100110011001100110", b"01000010110100110011001100110011"), -- 99.4 + 6.2 = 105.6
	(b"11000001011111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100000110011001100110011", b"00111111000110011001100110010000"), -- -15.8 + 16.4 = 0.599999
	(b"11000001100011000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010110110011001100110011", b"01000010000101010011001100110011"), -- -17.5 + 54.8 = 37.3
	(b"01000010010110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011101110011001100110011", b"11000000110111001100110011001000"), -- 54.9 + -61.8 = -6.9
	(b"11000010001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000100011001100110011", b"01000010010111100000000000000000"), -- -41.6 + 97.1 = 55.5
	(b"11000010100010101001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"11000010100100011001100110011010"), -- -69.3 + -3.5 = -72.8
	(b"01000010101111111001100110011010", b"00000000000000000000000000000000"),
	(b"11000000110110011001100110011010", b"01000010101100100000000000000000"), -- 95.8 + -6.8 = 89
	(b"01000001000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010010100000000000000000", b"11000010001001111001100110011010"), -- 8.6 + -50.5 = -41.9
	(b"11000001101111000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000001111001100110011010", b"01000001001001100110011001101000"), -- -23.5 + 33.9 = 10.4
	(b"11000010001000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111001100110011001100110", b"11000010001111100110011001100111"), -- -40.4 + -7.2 = -47.6
	(b"01000010011111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001111101110011001100110011", b"01000010101111001100110011001101"), -- 63.5 + 30.9 = 94.4
	(b"11000010011010101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111100001100110011001101", b"11000010101100011001100110011010"), -- -58.7 + -30.1 = -88.8
	(b"11000010010101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001000000000000000000", b"01000001111001001100110011001100"), -- -53.4 + 82 = 28.6
	(b"11000010100001110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101011000011001100110011", b"01000001100100110011001100110100"), -- -67.7 + 86.1 = 18.4
	(b"11000010100001110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010001100001100110011001101", b"11000010110111111100110011001100"), -- -67.7 + -44.2 = -111.9
	(b"01000010010111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111100001100110011001101", b"01000010101010111100110011001101"), -- 55.8 + 30.1 = 85.9
	(b"10111110100110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001110011100110011001100110", b"11000001110100001100110011001100"), -- -0.3 + -25.8 = -26.1
	(b"01000010100110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000010110011001100110", b"01000011001011100001100110011010"), -- 77.4 + 96.7 = 174.1
	(b"11000001111101001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111100110011001100110011010", b"11000001111010110011001100110011"), -- -30.6 + 1.2 = -29.4
	(b"11000001111011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110001010110011001100110", b"01000010100010011100110011001100"), -- -29.8 + 98.7 = 68.9
	(b"11000000111110011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001001011001100110011010", b"11000010010001001100110011001101"), -- -7.8 + -41.4 = -49.2
	(b"01000010100010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001011011100110011001100110", b"01000010101001011100110011001101"), -- 68 + 14.9 = 82.9
	(b"01000010001000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101001000011001100110011", b"11000010001010000000000000000000"), -- 40.1 + -82.1 = -42
	(b"01000010000001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011011010011001100110011", b"01000010101110001001100110011010"), -- 33 + 59.3 = 92.3
	(b"11000001110100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011011101100110011001101", b"01000010000001101100110011001101"), -- -26 + 59.7 = 33.7
	(b"11000010100110010110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001011100000000000000000", b"11000010000001001100110011001100"), -- -76.7 + 43.5 = -33.2
	(b"11000010011010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001011111001100110011001101", b"11000010001010011001100110011010"), -- -58.2 + 15.8 = -42.4
	(b"01000010010101000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001010011001100110011001101", b"01000010100000111001100110011010"), -- 53 + 12.8 = 65.8
	(b"01000010011100100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000101100000000000000000", b"01000010110001000000000000000000"), -- 60.5 + 37.5 = 98
	(b"01000010101001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000100011001100110011010", b"01000010111100000000000000000000"), -- 83.6 + 36.4 = 120
	(b"11000010101000011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011000101100110011001101", b"11000011000010011001100110011010"), -- -80.9 + -56.7 = -137.6
	(b"01000010100001110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010100011010110011001100110", b"01000011000010100011001100110011"), -- 67.5 + 70.7 = 138.2
	(b"11000010101100101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001010000000000000000000", b"11000010001111011001100110011010"), -- -89.4 + 42 = -47.4
	(b"11000001101100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111101001100110011001101", b"01000001000010000000000000000000"), -- -22.1 + 30.6 = 8.5
	(b"01000010000001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010001001111001100110011010", b"11000001000011100110011001101000"), -- 33 + -41.9 = -8.9
	(b"11000010001000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101001101100110011001101", b"11000010111110001001100110011010"), -- -40.9 + -83.4 = -124.3
	(b"11000010101101001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111110110011001100110011010", b"11000010101100010110011001100111"), -- -90.4 + 1.7 = -88.7
	(b"11000001111110001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101001010000000000000000", b"01000010010011011001100110011010"), -- -31.1 + 82.5 = 51.4
	(b"11000010000100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000000100010011001100110011010", b"11000010000000100110011001100111"), -- -36.9 + 4.3 = -32.6
	(b"01000001110110011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000111111001100110011010", b"01000010100001100011001100110100"), -- 27.2 + 39.9 = 67.1
	(b"01000000101010011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000011000000000000000000", b"01000010001000010011001100110011"), -- 5.3 + 35 = 40.3
	(b"11000010001000011001100110011010", b"00000000000000000000000000000000"),
	(b"10111111000000000000000000000000", b"11000010001000111001100110011010"), -- -40.4 + -0.5 = -40.9
	(b"11000010001111011001100110011010", b"00000000000000000000000000000000"),
	(b"11000001100011001100110011001101", b"11000010100000100000000000000000"), -- -47.4 + -17.6 = -65
	(b"11000010100110110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100101011100110011001101", b"11000011000110000110011001100110"), -- -77.5 + -74.9 = -152.4
	(b"11000001100110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010001010111001100110011010", b"01000001101111001100110011001110"), -- -19.3 + 42.9 = 23.6
	(b"11000010100100011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100010011001100110011010", b"11000011000011011001100110011010"), -- -72.8 + -68.8 = -141.6
	(b"11000001001101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011010111001100110011010", b"01000010001111100000000000000000"), -- -11.4 + 58.9 = 47.5
	(b"11000010100100101001100110011010", b"00000000000000000000000000000000"),
	(b"01000001101010000000000000000000", b"11000010010100010011001100110100"), -- -73.3 + 21 = -52.3
	(b"11000010110001001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101001001100110011001101", b"11000001011111100110011001101000"), -- -98.3 + 82.4 = -15.9
	(b"11000010100011000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000001100110011001101", b"01000001110100011001100110011100"), -- -70.2 + 96.4 = 26.2
	(b"11000010101101100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011010110011001100110", b"11000011001100011011001100110011"), -- -91 + -86.7 = -177.7
	(b"01000001011100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010101100110011001100110011", b"11000010100101001100110011001101"), -- 15.2 + -89.6 = -74.4
	(b"11000001110001110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111100110011001100110011", b"01000000101100000000000000000000"), -- -24.9 + 30.4 = 5.5
	(b"01000010101100000011001100110011", b"00000000000000000000000000000000"),
	(b"11000001111011100110011001100110", b"01000010011010010011001100110011"), -- 88.1 + -29.8 = 58.3
	(b"11000000100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010011000110011001100110", b"11000010010111011001100110011001"), -- -4.3 + -51.1 = -55.4
	(b"01000001100100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011001100000000000000000", b"01000010100101111001100110011010"), -- 18.3 + 57.5 = 75.8
	(b"11000010010000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011100110011001100110011", b"11000010010100001100110011001101"), -- -48.4 + -3.8 = -52.2
	(b"11000010011001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001000111001100110011010", b"11000001100010000000000000000000"), -- -57.9 + 40.9 = -17
	(b"11000010100001111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010100000000000000000", b"11000011000110001100110011001101"), -- -67.8 + -85 = -152.8
	(b"01000001001110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101000011001100110011", b"01000010101010111001100110011001"), -- 11.7 + 74.1 = 85.8
	(b"11000010010010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100101110000000000000000", b"01000001110010011001100110011010"), -- -50.3 + 75.5 = 25.2
	(b"11000010001010100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100001011001100110011010", b"11000001110011100110011001100110"), -- -42.5 + 16.7 = -25.8
	(b"11000001011001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010110000010000000000000000", b"01000010101001000110011001100110"), -- -14.3 + 96.5 = 82.2
	(b"01000001111010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100011001100110011010", b"01000001101000000000000000000000"), -- 29.1 + -9.1 = 20
	(b"01000010100010010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001110000000000000000", b"01000011000010000001100110011010"), -- 68.6 + 67.5 = 136.1
	(b"01000010101010000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011001100000000000000000", b"01000011000011011001100110011010"), -- 84.1 + 57.5 = 141.6
	(b"01000010010001000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000000000110011001100110", b"01000001100001110011001100110100"), -- 49 + -32.1 = 16.9
	(b"01000010010000000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100001010000000000000000", b"01000010111001010011001100110011"), -- 48.1 + 66.5 = 114.6
	(b"01000010101110000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101000011001100110011010", b"01000011001011010000000000000000"), -- 92.2 + 80.8 = 173
	(b"01000001100000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001011000110011001100110011", b"01000001111100100110011001100110"), -- 16.1 + 14.2 = 30.3
	(b"01000001000110000000000000000000", b"00000000000000000000000000000000"),
	(b"10111111110011001100110011001101", b"01000000111111001100110011001101"), -- 9.5 + -1.6 = 7.9
	(b"11000010010110000110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011101001100110011001101", b"01000000111000110011001100111000"), -- -54.1 + 61.2 = 7.1
	(b"11000010110001011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101100011100110011001101", b"11000001001000000000000000000000"), -- -98.9 + 88.9 = -10
	(b"01000010000111110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010000001101100110011001101", b"01000010100100110000000000000000"), -- 39.8 + 33.7 = 73.5
	(b"01000010011010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010110000101100110011001101", b"11000010000110100000000000000000"), -- 58.9 + -97.4 = -38.5
	(b"01000010001010010011001100110011", b"00000000000000000000000000000000"),
	(b"11000000110100000000000000000000", b"01000010000011110011001100110011"), -- 42.3 + -6.5 = 35.8
	(b"01000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001101000000000000000000", b"01000010010100000000000000000000"), -- 7 + 45 = 52
	(b"01000010101010110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010011011100110011001100110", b"01000011000100010100110011001100"), -- 85.7 + 59.6 = 145.3
	(b"11000010010111100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010011001000110011001100110", b"00111111110011001100110011000000"), -- -55.5 + 57.1 = 1.6
	(b"01000010101011110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000111100110011001101", b"11000001001001100110011001101000"), -- 87.5 + -97.9 = -10.4
	(b"01000010100010010000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000101100110011001100110", b"01000010011011000110011001100110"), -- 68.5 + -9.4 = 59.1
	(b"01000001010111100110011001100110", b"00000000000000000000000000000000"),
	(b"00111110110011001100110011001101", b"01000001011001001100110011001100"), -- 13.9 + 0.4 = 14.3
	(b"01000010101001011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001111011001100110011010", b"01000010000011011001100110011010"), -- 82.8 + -47.4 = 35.4
	(b"01000010001100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100011000000000000000000", b"11000001110100000000000000000000"), -- 44 + -70 = -26
	(b"01000010101001010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101011000110011001100110", b"11000000011011001100110011000000"), -- 82.5 + -86.2 = -3.7
	(b"11000010100010101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001111100000000000000000000", b"11000010110001101100110011001101"), -- -69.4 + -30 = -99.4
	(b"11000010010101101100110011001101", b"00000000000000000000000000000000"),
	(b"00111101110011001100110011001101", b"11000010010101100110011001100111"), -- -53.7 + 0.1 = -53.6
	(b"11000010011001111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000000000000000000000000", b"11000001110011110011001100110100"), -- -57.9 + 32 = -25.9
	(b"01000001110001001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101011001001100110011010", b"11000010011101101100110011001110"), -- 24.6 + -86.3 = -61.7
	(b"11000010101011000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000110001100110011001101", b"11000010111110000110011001100110"), -- -86 + -38.2 = -124.2
	(b"11000010010010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001001010110011001100110011", b"11000010011101100000000000000000"), -- -50.8 + -10.7 = -61.5
	(b"01000010000010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111110100110011001100110", b"01000000001011001100110011010000"), -- 34 + -31.3 = 2.7
	(b"01000010101010111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011011000000000000000000", b"01000001110101100110011001101000"), -- 85.8 + -59 = 26.8
	(b"11000010010100100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001110010000000000000000000", b"11000001110111001100110011001100"), -- -52.6 + 25 = -27.6
	(b"11000001110001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010000101110011001100110011", b"11000010011110100110011001100110"), -- -24.8 + -37.8 = -62.6
	(b"11000001000110110011001100110011", b"00000000000000000000000000000000"),
	(b"11000000111111001100110011001101", b"11000001100011001100110011001101"), -- -9.7 + -7.9 = -17.6
	(b"11000010101110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001000110000000000000000000", b"11000010101001111100110011001101"), -- -93.4 + 9.5 = -83.9
	(b"01000001111100100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001001000110011001100110011", b"01000001101000001100110011001100"), -- 30.3 + -10.2 = 20.1
	(b"01000010100011110000000000000000", b"00000000000000000000000000000000"),
	(b"01000001000101100110011001100110", b"01000010101000011100110011001101"), -- 71.5 + 9.4 = 80.9
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011010111001100110011010", b"11000010100000011100110011001101"), -- -6 + -58.9 = -64.9
	(b"11000010100110010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100101011100110011001101", b"11000011000101111001100110011010"), -- -76.7 + -74.9 = -151.6
	(b"11000001001100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000010110011001100110011", b"11000010001101110011001100110011"), -- -11 + -34.8 = -45.8
	(b"11000000111000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001111111001100110011001101", b"11000010000110100110011001100110"), -- -7 + -31.6 = -38.6
	(b"01000001011010000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101000111100110011001101", b"01000010110000001100110011001101"), -- 14.5 + 81.9 = 96.4
	(b"01000000000011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000001000100000000000000000000", b"11000000110110011001100110011010"), -- 2.2 + -9 = -6.8
	(b"11000010101001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101001011001100110011010", b"11000010011101010011001100110011"), -- -82 + 20.7 = -61.3
	(b"11000010100111110110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101110000000000000000000", b"11000011001010111011001100110011"), -- -79.7 + -92 = -171.7
	(b"01000010101110010011001100110011", b"00000000000000000000000000000000"),
	(b"01000001011001001100110011001101", b"01000010110101011100110011001101"), -- 92.6 + 14.3 = 106.9
	(b"11000010100000000110011001100110", b"00000000000000000000000000000000"),
	(b"11000000000110011001100110011010", b"11000010100001010011001100110011"), -- -64.2 + -2.4 = -66.6
	(b"11000001111101110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001001101100110011001101", b"01000001001011001100110011001110"), -- -30.9 + 41.7 = 10.8
	(b"11000010101011000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100001100011001100110011", b"11000011000110010100110011001100"), -- -86.2 + -67.1 = -153.3
	(b"01000010000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001100101110011001100110011", b"01000001100001011001100110011001"), -- 35.6 + -18.9 = 16.7
	(b"11000010100100010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100100111100110011001101", b"11000011000100100110011001100110"), -- -72.5 + -73.9 = -146.4
	(b"01000010100111110000000000000000", b"00000000000000000000000000000000"),
	(b"01000010001011000000000000000000", b"01000010111101010000000000000000"), -- 79.5 + 43 = 122.5
	(b"01000010101111010110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001111100110011001101", b"11000000101001100110011001110000"), -- 94.7 + -99.9 = -5.2
	(b"01000010001010000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110000101001100110011010", b"11000010010111001100110011001110"), -- 42.1 + -97.3 = -55.2
	(b"01000010010101010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001101100110011001101", b"01000010111100010110011001100110"), -- 53.3 + 67.4 = 120.7
	(b"01000010100100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000000110011001100110", b"11000001110000011001100110011000"), -- 72 + -96.2 = -24.2
	(b"11000000110000000000000000000000", b"00000000000000000000000000000000"),
	(b"01000001101100100110011001100110", b"01000001100000100110011001100110"), -- -6 + 22.3 = 16.3
	(b"11000010010100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010000001000000000000000000", b"11000001100110110011001100110100"), -- -52.4 + 33 = -19.4
	(b"01000001110000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"01000001111000000000000000000000"), -- 24.4 + 3.6 = 28
	(b"01000001100010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111110011001100110011010", b"01000001000101100110011001100111"), -- 17.2 + -7.8 = 9.4
	(b"01000010000010000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110000101001100110011010", b"11000010011111001100110011001110"), -- 34.1 + -97.3 = -63.2
	(b"01000010100000110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011100111001100110011010", b"01000010111111010000000000000000"), -- 65.6 + 60.9 = 126.5
	(b"10111111000000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010100101111001100110011010", b"11000010100110001001100110011010"), -- -0.5 + -75.8 = -76.3
	(b"11000001111101011001100110011010", b"00000000000000000000000000000000"),
	(b"11000000111100110011001100110011", b"11000010000110010011001100110011"), -- -30.7 + -7.6 = -38.3
	(b"01000010001001000110011001100110", b"00000000000000000000000000000000"),
	(b"01000001011000011001100110011010", b"01000010010111001100110011001100"), -- 41.1 + 14.1 = 55.2
	(b"11000010101000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000010110011001100110", b"10111101110011001101000000000000"), -- -80.8 + 80.7 = -0.100006
	(b"01000010100010111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101100000011001100110011", b"01000011000111100000000000000000"), -- 69.9 + 88.1 = 158
	(b"11000000100101100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000011001100110011001100110", b"10111111100011001100110011001100"), -- -4.7 + 3.6 = -1.1
	(b"11000010100111011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010001001000110011001100110", b"11000010111100000000000000000000"), -- -78.9 + -41.1 = -120
	(b"11000010010011110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010000100100000000000000000", b"11000010101100001001100110011010"), -- -51.8 + -36.5 = -88.3
	(b"01000001100010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101111001100110011001101", b"01000010001001000000000000000000"), -- 17.4 + 23.6 = 41
	(b"11000010100001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010101110011001100110011", b"11000010111100101100110011001100"), -- -67.6 + -53.8 = -121.4
	(b"11000010101001100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010010110011001100110011010", b"11000001111001001100110011001100"), -- -83 + 54.4 = -28.6
	(b"11000010010000100000000000000000", b"00000000000000000000000000000000"),
	(b"01000000010000000000000000000000", b"11000010001101100000000000000000"), -- -48.5 + 3 = -45.5
	(b"11000001101011011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101111000110011001100110", b"11000010111001111100110011001100"), -- -21.7 + -94.2 = -115.9
	(b"01000010101000110000000000000000", b"00000000000000000000000000000000"),
	(b"01000000100110011001100110011010", b"01000010101011001001100110011010"), -- 81.5 + 4.8 = 86.3
	(b"11000001101001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000000010100110011001100110011", b"11000001100011000000000000000000"), -- -20.8 + 3.3 = -17.5
	(b"01000010101000111001100110011010", b"00000000000000000000000000000000"),
	(b"11000000011000000000000000000000", b"01000010100111001001100110011010"), -- 81.8 + -3.5 = 78.3
	(b"01000010100101110000000000000000", b"00000000000000000000000000000000"),
	(b"01000000000011001100110011001101", b"01000010100110110110011001100110"), -- 75.5 + 2.2 = 77.7
	(b"11000010010111001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010000011000000000000000000", b"11000010101101000110011001100110"), -- -55.2 + -35 = -90.2
	(b"11000010100001010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100011110011001100110011", b"01000000101000000000000000000000"), -- -66.6 + 71.6 = 5
	(b"01000010001100111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010100110110011001100110011", b"11000010000000101100110011001100"), -- 44.9 + -77.6 = -32.7
	(b"01000010001100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001011010000000000000000000", b"01000010011010111001100110011010"), -- 44.4 + 14.5 = 58.9
	(b"11000010000011111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101000111001100110011010", b"01000010001101111001100110011010"), -- -35.9 + 81.8 = 45.9
	(b"11000010001101001100110011001101", b"00000000000000000000000000000000"),
	(b"01000001111111000000000000000000", b"11000001010110110011001100110100"), -- -45.2 + 31.5 = -13.7
	(b"01000001111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001001010011001100110011010", b"01000001100110110011001100110011"), -- 30 + -10.6 = 19.4
	(b"01000010010011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101100000110011001100110", b"11000010000100101100110011001100"), -- 51.5 + -88.2 = -36.7
	(b"01000010100010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010010010001100110011001101", b"01000001100100011001100110011010"), -- 68.4 + -50.2 = 18.2
	(b"11000010011010110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100100110000000000000000", b"11000011000001000100110011001101"), -- -58.8 + -73.5 = -132.3
	(b"11000010101001000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101010010000000000000000", b"01000000001000000000000000000000"), -- -82 + 84.5 = 2.5
	(b"11000000100001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001010011001100110011001101", b"11000001100010000000000000000000"), -- -4.2 + -12.8 = -17
	(b"11000010101100010000000000000000", b"00000000000000000000000000000000"),
	(b"11000010010011100000000000000000", b"11000011000011000000000000000000"), -- -88.5 + -51.5 = -140
	(b"01000001010100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001111011100110011001100110", b"01000010001011000000000000000000"), -- 13.2 + 29.8 = 43
	(b"01000010101110110000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011111010011001100110011", b"01000001111100011001100110011010"), -- 93.5 + -63.3 = 30.2
	(b"11000010001110100000000000000000", b"00000000000000000000000000000000"),
	(b"00111111000110011001100110011010", b"11000010001101111001100110011010"), -- -46.5 + 0.6 = -45.9
	(b"11000000111100000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010101110101001100110011010", b"11000010110010011001100110011010"), -- -7.5 + -93.3 = -100.8
	(b"01000010101010001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100010011100110011001101", b"01000011000110010100110011001101"), -- 84.4 + 68.9 = 153.3
	(b"01000010101000010110011001100110", b"00000000000000000000000000000000"),
	(b"11000001000110000000000000000000", b"01000010100011100110011001100110"), -- 80.7 + -9.5 = 71.2
	(b"01000001101101000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011010111001100110011010", b"11000010000100011001100110011010"), -- 22.5 + -58.9 = -36.4
	(b"11000010011011100000000000000000", b"00000000000000000000000000000000"),
	(b"01000010000000110011001100110011", b"11000001110101011001100110011010"), -- -59.5 + 32.8 = -26.7
	(b"11000010010101000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010110001100011001100110011", b"11000011000110000011001100110011"), -- -53.1 + -99.1 = -152.2
	(b"11000010100110000011001100110011", b"00000000000000000000000000000000"),
	(b"01000010011110101100110011001101", b"11000001010101100110011001100100"), -- -76.1 + 62.7 = -13.4
	(b"11000001010011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101001011001100110011010", b"11000010000001100110011001100110"), -- -12.9 + -20.7 = -33.6
	(b"11000001011110110011001100110011", b"00000000000000000000000000000000"),
	(b"01000001101111000000000000000000", b"01000000111110011001100110011010"), -- -15.7 + 23.5 = 7.8
	(b"11000010001011010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001001000011001100110011010", b"11000010010101011001100110011010"), -- -43.3 + -10.1 = -53.4
	(b"01000010100110100110011001100110", b"00000000000000000000000000000000"),
	(b"01000001101011001100110011001101", b"01000010110001011001100110011001"), -- 77.2 + 21.6 = 98.8
	(b"11000010101010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101111111100110011001101", b"11000011001101000100110011001101"), -- -84.4 + -95.9 = -180.3
	(b"11000010100011100000000000000000", b"00000000000000000000000000000000"),
	(b"11000001110001000000000000000000", b"11000010101111110000000000000000"), -- -71 + -24.5 = -95.5
	(b"11000010100011101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010101010110000000000000000", b"01000001011000110011001100110000"), -- -71.3 + 85.5 = 14.2
	(b"11000010010111100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010110000100110011001100110", b"01000010001001100110011001100110"), -- -55.6 + 97.2 = 41.6
	(b"11000001100001001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001101100110011001100110", b"01000001111001111111111111111111"), -- -16.6 + 45.6 = 29
	(b"11000010001010101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101001100110011001100110", b"01000010001000011111111111111111"), -- -42.7 + 83.2 = 40.5
	(b"01000010000011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010100100000110011001100110", b"11000010000100100110011001100110"), -- 35.6 + -72.2 = -36.6
	(b"11000010100100011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100111011001100110011010", b"11000010010101000110011001100111"), -- -72.8 + 19.7 = -53.1
	(b"01000010100010001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010001110111001100110011010", b"01000001101010110011001100110100"), -- 68.3 + -46.9 = 21.4
	(b"11000010100001101001100110011010", b"00000000000000000000000000000000"),
	(b"10111111001100110011001100110011", b"11000010100010000000000000000000"), -- -67.3 + -0.7 = -68
	(b"11000000110000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010001101010011001100110011", b"11000010010011011001100110011001"), -- -6.1 + -45.3 = -51.4
	(b"11000001010010110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110101100110011001101", b"01000010100000010110011001100111"), -- -12.7 + 77.4 = 64.7
	(b"01000000001001100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010010010100000000000000000", b"01000010010101000110011001100110"), -- 2.6 + 50.5 = 53.1
	(b"01000010010111101100110011001101", b"00000000000000000000000000000000"),
	(b"11000001110101000000000000000000", b"01000001111010011001100110011010"), -- 55.7 + -26.5 = 29.2
	(b"11000001100000011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010011110110011001100110011", b"11000010100111100000000000000000"), -- -16.2 + -62.8 = -79
	(b"11000010100111011001100110011010", b"00000000000000000000000000000000"),
	(b"01000001100100011001100110011010", b"11000010011100100110011001100111"), -- -78.8 + 18.2 = -60.6
	(b"01000001110111001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101000110110011001100110", b"01000010110110101001100110011001"), -- 27.6 + 81.7 = 109.3
	(b"11000010010111010011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100001100011001100110011", b"01000001001111001100110011001100"), -- -55.3 + 67.1 = 11.8
	(b"00111111111001100110011001100110", b"00000000000000000000000000000000"),
	(b"11000010101101001100110011001101", b"11000010101100010011001100110011"), -- 1.8 + -90.4 = -88.6
	(b"01000001110000100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101000011001100110011010", b"01000000100000110011001100110000"), -- 24.3 + -20.2 = 4.1
	(b"11000010100011000110011001100110", b"00000000000000000000000000000000"),
	(b"11000010010001011001100110011010", b"11000010111011110011001100110011"), -- -70.2 + -49.4 = -119.6
	(b"11000001101000001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010010001100110011001100110", b"01000001111010111111111111111111"), -- -20.1 + 49.6 = 29.5
	(b"01000010011100001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010100110010000000000000000", b"01000011000010001011001100110011"), -- 60.2 + 76.5 = 136.7
	(b"11000010100111001001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101000001100110011001101", b"11000011000111101011001100110100"), -- -78.3 + -80.4 = -158.7
	(b"01000001010100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010010110001100110011001101", b"11000010001001000000000000000000"), -- 13.2 + -54.2 = -41
	(b"01000010000110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011100100110011001100110", b"11000001101100100110011001100110"), -- 38.3 + -60.6 = -22.3
	(b"11000010000000101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100000011001100110011010", b"11000001100001000000000000000000"), -- -32.7 + 16.2 = -16.5
	(b"11000010001100100000000000000000", b"00000000000000000000000000000000"),
	(b"11000010011000001100110011001101", b"11000010110010010110011001100110"), -- -44.5 + -56.2 = -100.7
	(b"01000010010101010011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110110011001100110011010", b"01000010011100000110011001100110"), -- 53.3 + 6.8 = 60.1
	(b"11000010101010011100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101111000000000000000000", b"11000011001100101110011001100110"), -- -84.9 + -94 = -178.9
	(b"11000010110001001001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010011001100110011001101", b"11000010001111000110011001100111"), -- -98.3 + 51.2 = -47.1
	(b"11000010101001110011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101001000000000000000000", b"11000010110100000011001100110011"), -- -83.6 + -20.5 = -104.1
	(b"11000010000010011001100110011010", b"00000000000000000000000000000000"),
	(b"11000010101010111001100110011010", b"11000010111100000110011001100111"), -- -34.4 + -85.8 = -120.2
	(b"01000010010110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100101001100110011001101", b"11000001101000001100110011001110"), -- 54.3 + -74.4 = -20.1
	(b"01000010010101111001100110011010", b"00000000000000000000000000000000"),
	(b"01000001110011011001100110011010", b"01000010100111110011001100110100"), -- 53.9 + 25.7 = 79.6
	(b"11000010100101011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100010110011001100110011", b"11000000101001100110011001110000"), -- -74.8 + 69.6 = -5.2
	(b"01000010010000110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011101000110011001100110", b"11000001010001001100110011001100"), -- 48.8 + -61.1 = -12.3
	(b"01000010101001110110011001100110", b"00000000000000000000000000000000"),
	(b"01000010101111110000000000000000", b"01000011001100110011001100110011"), -- 83.7 + 95.5 = 179.2
	(b"01000010100110011100110011001101", b"00000000000000000000000000000000"),
	(b"01000010101110001100110011001101", b"01000011001010010100110011001101"), -- 76.9 + 92.4 = 169.3
	(b"01000010011010000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001101010110011001100110011", b"01000010000100100110011001100110"), -- 58 + -21.4 = 36.6
	(b"01000001101100001100110011001101", b"00000000000000000000000000000000"),
	(b"00111111000000000000000000000000", b"01000001101101001100110011001101"), -- 22.1 + 0.5 = 22.6
	(b"11000010100110111001100110011010", b"00000000000000000000000000000000"),
	(b"11000010010000000110011001100110", b"11000010111110111100110011001101"), -- -77.8 + -48.1 = -125.9
	(b"11000000101100000000000000000000", b"00000000000000000000000000000000"),
	(b"01000010101000100011001100110011", b"01000010100101110011001100110011"), -- -5.5 + 81.1 = 75.6
	(b"11000010101110000011001100110011", b"00000000000000000000000000000000"),
	(b"11000000101111001100110011001101", b"11000010110001000000000000000000"), -- -92.1 + -5.9 = -98
	(b"01000010101010001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010101000110110011001100110", b"01000000001011001100110011100000"), -- 84.4 + -81.7 = 2.7
	(b"11000010101000011001100110011010", b"00000000000000000000000000000000"),
	(b"01000010001001011001100110011010", b"11000010000111011001100110011010"), -- -80.8 + 41.4 = -39.4
	(b"11000010000011111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100001010110011001100110", b"01000001111101100110011001100100"), -- -35.9 + 66.7 = 30.8
	(b"11000001100000001100110011001101", b"00000000000000000000000000000000"),
	(b"11000010011101111001100110011010", b"11000010100111000000000000000000"), -- -16.1 + -61.9 = -78
	(b"11000000101100110011001100110011", b"00000000000000000000000000000000"),
	(b"11000010100110100000000000000000", b"11000010101001010011001100110011"), -- -5.6 + -77 = -82.6
	(b"01000010010110101100110011001101", b"00000000000000000000000000000000"),
	(b"01000001110010001100110011001101", b"01000010100111111001100110011010"), -- 54.7 + 25.1 = 79.8
	(b"01000010100010010011001100110011", b"00000000000000000000000000000000"),
	(b"11000001101000110011001100110011", b"01000010010000001100110011001100"), -- 68.6 + -20.4 = 48.2
	(b"01000010100000100000000000000000", b"00000000000000000000000000000000"),
	(b"01000001100001110011001100110011", b"01000010101000111100110011001101"), -- 65 + 16.9 = 81.9
	(b"01000010100110000000000000000000", b"00000000000000000000000000000000"),
	(b"11000001000100110011001100110011", b"01000010100001011001100110011010"), -- 76 + -9.2 = 66.8
	(b"11000001001011100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001011011100110011001100110", b"11000001110011100110011001100110"), -- -10.9 + -14.9 = -25.8
	(b"11000010100100111001100110011010", b"00000000000000000000000000000000"),
	(b"01000010100010000011001100110011", b"11000000101101100110011001110000"), -- -73.8 + 68.1 = -5.7
	(b"01000010100101111100110011001101", b"00000000000000000000000000000000"),
	(b"01000001100001011001100110011010", b"01000010101110010011001100110100"), -- 75.9 + 16.7 = 92.6
	(b"00111111010011001100110011001101", b"00000000000000000000000000000000"),
	(b"11000000100010011001100110011010", b"11000000011000000000000000000001"), -- 0.8 + -4.3 = -3.5
	(b"01000010110000110110011001100110", b"00000000000000000000000000000000"),
	(b"11000001101001100110011001100110", b"01000010100110011100110011001100"), -- 97.7 + -20.8 = 76.9
	(b"01000001011000000000000000000000", b"00000000000000000000000000000000"),
	(b"11000010000000000000000000000000", b"11000001100100000000000000000000"), -- 14 + -32 = -18
	(b"01000010000110010011001100110011", b"00000000000000000000000000000000"),
	(b"11000010011011101100110011001101", b"11000001101010110011001100110100"), -- 38.3 + -59.7 = -21.4
	(b"11000000101011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010001000111001100110011010", b"01000010000011100000000000000000"), -- -5.4 + 40.9 = 35.5
	(b"11000010001011110011001100110011", b"00000000000000000000000000000000"),
	(b"01000010100110110110011001100110", b"01000010000001111001100110011001"), -- -43.8 + 77.7 = 33.9
	(b"01000000001100110011001100110011", b"00000000000000000000000000000000"),
	(b"01000000110000000000000000000000", b"01000001000011001100110011001101"), -- 2.8 + 6 = 8.8
	(b"11000010011011001100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000011111001100110011010", b"11000001101110100110011001100110"), -- -59.2 + 35.9 = -23.3
	(b"01000010100011100110011001100110", b"00000000000000000000000000000000"),
	(b"01000010100010001100110011001101", b"01000011000010111001100110011010"), -- 71.2 + 68.4 = 139.6
	(b"11000010101110111100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000101001100110011001101", b"11000010011000101100110011001101"), -- -93.9 + 37.2 = -56.7
	(b"11000010011100101100110011001101", b"00000000000000000000000000000000"),
	(b"01000010000101010011001100110011", b"11000001101110110011001100110100"), -- -60.7 + 37.3 = -23.4
	(b"01000010101110101001100110011010", b"00000000000000000000000000000000"),
	(b"01000010010001001100110011001101", b"01000011000011101000000000000000"), -- 93.3 + 49.2 = 142.5
	(b"01000010100101100110011001100110", b"00000000000000000000000000000000"),
	(b"11000001110100110011001100110011", b"01000010010000110011001100110010"), -- 75.2 + -26.4 = 48.8
	(b"01000010100010100011001100110011", b"00000000000000000000000000000000"),
	(b"01000010001000110011001100110011", b"01000010110110111100110011001100"), -- 69.1 + 40.8 = 109.9

	(b"01000010100111111011010111100000", b"00000000000000000000000000000000"),
	(b"11000010101011010010000001101101", b"11000000110101101010100011010000"), -- 79.8552 + -86.5633 = -6.70811
	(b"01000010100111010100011011000001", b"00000000000000000000000000000000"),
	(b"11000001000000111111011001010000", b"01000010100011001100011111110111"), -- 78.6382 + -8.24763 = 70.3906
	(b"11000001111101001010011000111000", b"00000000000000000000000000000000"),
	(b"01000010110000011111101010011100", b"01000010100001001101000100001110"), -- -30.5812 + 96.9895 = 66.4083
	(b"11000010101110111011010000110010", b"00000000000000000000000000000000"),
	(b"11000001101010110100110111110000", b"11000010111001101000011110101110"), -- -93.8519 + -21.4131 = -115.265
	(b"11000001100111100101011011010000", b"00000000000000000000000000000000"),
	(b"11000010010111101001010001011010", b"11000010100101101101111111100001"), -- -19.7924 + -55.6449 = -75.4373
	(b"11000001100111110101100010001000", b"00000000000000000000000000000000"),
	(b"01000001100101110111000111110000", b"10111111011111001101001100000000"), -- -19.9182 + 18.9306 = -0.987595
	(b"11000000101111100101111101110000", b"00000000000000000000000000000000"),
	(b"01000001101001011100011100110000", b"01000001011011000101111010101000"), -- -5.94915 + 20.7223 = 14.7731
	(b"11000010100110000111101101000110", b"00000000000000000000000000000000"),
	(b"11000010010010001000000100000110", b"11000010111111001011101111001001"), -- -76.2408 + -50.126 = -126.367
	(b"01000010001101011000001111110000", b"00000000000000000000000000000000"),
	(b"11000010010010001001101001001001", b"11000000100110001011001011001000"), -- 45.3788 + -50.1507 = -4.77182
	(b"11000010100011001100101101111110", b"00000000000000000000000000000000"),
	(b"11000000011100011000101111000000", b"11000010100101000101011111011100"), -- -70.3974 + -3.77415 = -74.1716
	(b"01000010110001000010100111011101", b"00000000000000000000000000000000"),
	(b"01000010011111000101011011101100", b"01000011001000010010101010101010"), -- 98.0818 + 63.0849 = 161.167
	(b"11000000101011010011000101100000", b"00000000000000000000000000000000"),
	(b"11000010101011011100011000111100", b"11000010101110001001100101010010"), -- -5.41228 + -86.8872 = -92.2995
	(b"11000010101110110110011100010100", b"00000000000000000000000000000000"),
	(b"01000010001101101100000101001010", b"11000010010000000000110011011110"), -- -93.7013 + 45.6888 = -48.0126
	(b"11000010001010110001100101001100", b"00000000000000000000000000000000"),
	(b"01000010101111011110101010101000", b"01000010010100001011110000000100"), -- -42.7747 + 94.9583 = 52.1836
	(b"11000010011000110001001111001100", b"00000000000000000000000000000000"),
	(b"11000001100111011110000110001100", b"11000010100110010000001001001001"), -- -56.7693 + -19.7351 = -76.5045
	(b"01000001111001110100000011110100", b"00000000000000000000000000000000"),
	(b"01000001001110110001000111000000", b"01000010001000100110010011101010"), -- 28.9067 + 11.6918 = 40.5985
	(b"11000010101000110101110011000110", b"00000000000000000000000000000000"),
	(b"01000010100001011110000101110110", b"11000001011010111101101010000000"), -- -81.6812 + 66.9404 = -14.7408
	(b"11000010100111010010110011100110", b"00000000000000000000000000000000"),
	(b"01000010100111101000110111101111", b"00111111001100001000010010000000"), -- -78.5877 + 79.2772 = 0.689522
	(b"01000000100000100111111001010000", b"00000000000000000000000000000000"),
	(b"11000000101000110101011111110000", b"10111111100000110110011010000000"), -- 4.07792 + -5.10448 = -1.02657
	(b"01000010101011010111101000100101", b"00000000000000000000000000000000"),
	(b"11000010101000100010011110000010", b"01000000101101010010101000110000"), -- 86.7386 + -81.0772 = 5.6614
	(b"11000001100111001001101111000000", b"00000000000000000000000000000000"),
	(b"11000010100010110110011011001100", b"11000010101100101000110110111100"), -- -19.576 + -69.7008 = -89.2768
	(b"01000001101011100100101001100000", b"00000000000000000000000000000000"),
	(b"01000010100001010011011100010100", b"01000010101100001100100110101100"), -- 21.7863 + 66.6076 = 88.3939
	(b"11000010001011010111000010011000", b"00000000000000000000000000000000"),
	(b"01000010101111010110010110111010", b"01000010010011010101101011011100"), -- -43.36 + 94.6987 = 51.3387
	(b"01000010100000010100100100111000", b"00000000000000000000000000000000"),
	(b"11000010100110101011111001010010", b"11000001010010111010100011010000"), -- 64.643 + -77.3717 = -12.7287
	(b"11000010000111101110111110000101", b"00000000000000000000000000000000"),
	(b"01000010010011000000001011001011", b"01000001001101000100110100011000"), -- -39.7339 + 51.0027 = 11.2688
	(b"11000010101011010111000110100010", b"00000000000000000000000000000000"),
	(b"01000001000110001000011000001000", b"11000010100110100110000011100001"), -- -86.7219 + 9.53272 = -77.1892
	(b"11000001110110001101000101100000", b"00000000000000000000000000000000"),
	(b"01000010101111111101111100100010", b"01000010100010011010101011001010"), -- -27.1022 + 95.9358 = 68.8336
	(b"11000001100100100000001011100000", b"00000000000000000000000000000000"),
	(b"01000010100111111010000011010100", b"01000010011101100100000000111000"), -- -18.2514 + 79.8141 = 61.5627
	(b"01000001111110011110110110001000", b"00000000000000000000000000000000"),
	(b"01000010011111000010001001101100", b"01000010101111001000110010011000"), -- 31.241 + 63.0336 = 94.2746
	(b"11000010001101011010010010110010", b"00000000000000000000000000000000"),
	(b"11000010001000100000000110001000", b"11000010101010111101001100011101"), -- -45.4108 + -40.5015 = -85.9123
	(b"11000001101011011110101000111100", b"00000000000000000000000000000000"),
	(b"11000010010110101010101100010000", b"11000010100110001101000000010111"), -- -21.7394 + -54.6671 = -76.4064
	(b"11000010011111110100000000111000", b"00000000000000000000000000000000"),
	(b"11000010001100111011101011111001", b"11000010110110010111110110011000"), -- -63.8127 + -44.9326 = -108.745
	(b"01000001110110100001101001100000", b"00000000000000000000000000000000"),
	(b"01000010011100000001000010001100", b"01000010101011101000111011011110"), -- 27.2629 + 60.0162 = 87.279
	(b"01000010001110101100111111010100", b"00000000000000000000000000000000"),
	(b"01000010101000000110010000111010", b"01000010111111011100110000100100"), -- 46.703 + 80.1958 = 126.899
	(b"01000010101110010000010111101100", b"00000000000000000000000000000000"),
	(b"01000010100011010001011011000100", b"01000011001000110000111001011000"), -- 92.5116 + 70.5445 = 163.056
	(b"01000010100100011100000000010000", b"00000000000000000000000000000000"),
	(b"11000010100000100101000010010110", b"01000000111101101111011110100000"), -- 72.8751 + -65.1574 = 7.71773
	(b"11000010010001001011100010100101", b"00000000000000000000000000000000"),
	(b"11000010100100110010000000000100", b"11000010111101010111110001010110"), -- -49.1803 + -73.5625 = -122.743
	(b"01000001100001100010001000101000", b"00000000000000000000000000000000"),
	(b"11000010100010110010110110000000", b"11000010010100110100100111101100"), -- 16.7667 + -69.5889 = -52.8222
	(b"01000010000000001111001011100000", b"00000000000000000000000000000000"),
	(b"11000001011110100010000011100000", b"01000001100001001101010101010000"), -- 32.2372 + -15.633 = 16.6042
	(b"11000010000011101001101111000000", b"00000000000000000000000000000000"),
	(b"11000001100100011100000011110000", b"11000010010101110111110000111000"), -- -35.6521 + -18.2192 = -53.8713
	(b"01000000111000011010011110110000", b"00000000000000000000000000000000"),
	(b"11000010011001001000010100011000", b"11000010010010000101000000100010"), -- 7.05172 + -57.13 = -50.0783
	(b"01000001001011011011011000111000", b"00000000000000000000000000000000"),
	(b"11000010101111110101100011111000", b"11000010101010011010001000110001"), -- 10.857 + -95.6738 = -84.8168
	(b"01000010001100111111010001100100", b"00000000000000000000000000000000"),
	(b"00111110010111100011111000000000", b"01000010001101001101001010100010"), -- 44.9887 + 0.217033 = 45.2057
	(b"11000001010110010100100100111000", b"00000000000000000000000000000000"),
	(b"01000010010100001000011101011010", b"01000010000110100011010100001100"), -- -13.5804 + 52.1322 = 38.5518
	(b"11000010101110000011001011110110", b"00000000000000000000000000000000"),
	(b"01000010001001010111011110000100", b"11000010010010101110111001101000"), -- -92.0995 + 41.3667 = -50.7328
	(b"11000010011110001001011001101001", b"00000000000000000000000000000000"),
	(b"01000001010100110101111011011000", b"11000010010000111011111010110011"), -- -62.1469 + 13.2107 = -48.9362
	(b"11000010101011111010000011101011", b"00000000000000000000000000000000"),
	(b"11000001000011000110101111010000", b"11000010110000010010111001100101"), -- -87.8143 + -8.77632 = -96.5906
	(b"01000010110001011011010000100010", b"00000000000000000000000000000000"),
	(b"11000010000110010010001111110001", b"01000010011100100100010001010011"), -- 98.8518 + -38.2851 = 60.5667
	(b"11000010100001100011111110001110", b"00000000000000000000000000000000"),
	(b"01000010110000110010110010001110", b"01000001111100111011010000000000"), -- -67.1241 + 97.587 = 30.4629
	(b"01000010101100111111001001110101", b"00000000000000000000000000000000"),
	(b"10111110001001101001110000000000", b"01000010101100111001111100100111"), -- 89.9735 + -0.162704 = 89.8108
	(b"01000010001010111000110110000000", b"00000000000000000000000000000000"),
	(b"11000010101110101000111010000110", b"11000010010010011000111110001100"), -- 42.8882 + -93.2784 = -50.3902
	(b"11000010000101100010010001101000", b"00000000000000000000000000000000"),
	(b"11000010100110111111000000010011", b"11000010111001110000001001000111"), -- -37.5356 + -77.9689 = -115.504
	(b"11000010100100111101100010011000", b"00000000000000000000000000000000"),
	(b"01000001100111100110111110110000", b"11000010010110000111100101011000"), -- -73.923 + 19.8045 = -54.1185
	(b"01000010010101110110000110010100", b"00000000000000000000000000000000"),
	(b"11000010101000001110011101110001", b"11000001110101001101101010011100"), -- 53.8453 + -80.452 = -26.6067
	(b"00111111110000100100110001000000", b"00000000000000000000000000000000"),
	(b"01000010001010000111001100011100", b"01000010001011101000010101111110"), -- 1.51795 + 42.1124 = 43.6304
	(b"11000010100001100010000100101110", b"00000000000000000000000000000000"),
	(b"01000010011100011100001000111110", b"11000000110101000000000011110000"), -- -67.0648 + 60.4397 = -6.62511
	(b"01000010100001100100110110101000", b"00000000000000000000000000000000"),
	(b"01000000011100010110000110000000", b"01000010100011011101100010110100"), -- 67.1517 + 3.77158 = 70.9232
	(b"11000010100011101011000101111101", b"00000000000000000000000000000000"),
	(b"11000010010011010010011100101111", b"11000010111101010100010100010100"), -- -71.3467 + -51.2883 = -122.635
	(b"01000010101001110011010000000000", b"00000000000000000000000000000000"),
	(b"11000010010001011101001000011100", b"01000010000010001001010111100100"), -- 83.6016 + -49.4552 = 34.1464
	(b"11000010100111100110000101011011", b"00000000000000000000000000000000"),
	(b"01000010100010001110001100100010", b"11000001001010111111000111001000"), -- -79.1901 + 68.4436 = -10.7465
	(b"11000010010001111010001010010000", b"00000000000000000000000000000000"),
	(b"11000000000101011111010110100000", b"11000010010100010000000111101010"), -- -49.9088 + -2.34312 = -52.2519
	(b"11000010011001000110001000010010", b"00000000000000000000000000000000"),
	(b"01000010011011001001001000000000", b"01000000000000101111111011100000"), -- -57.0958 + 59.1426 = 2.04681
	(b"01000000101000101101110000000000", b"00000000000000000000000000000000"),
	(b"11000010100011100001100110111000", b"11000010100000111110101111111000"), -- 5.08936 + -71.0502 = -65.9609
	(b"11000001001101100110000011001000", b"00000000000000000000000000000000"),
	(b"01000010010010111001011110001110", b"01000010000111011111111101011100"), -- -11.3986 + 50.898 = 39.4994
	(b"11000010000110110110111100101101", b"00000000000000000000000000000000"),
	(b"01000010110001001000000100100100", b"01000010011011011001001100011011"), -- -38.8586 + 98.2522 = 59.3937
	(b"11000010011001110111111010000100", b"00000000000000000000000000000000"),
	(b"11000010100000011110001100101010", b"11000010111101011010001001101100"), -- -57.8736 + -64.9437 = -122.817
	(b"11000010000010111110111101110100", b"00000000000000000000000000000000"),
	(b"01000010001001100010000100100011", b"01000000110100011000110101111000"), -- -34.9838 + 41.5324 = 6.54852
	(b"11000010100000010000111100011010", b"00000000000000000000000000000000"),
	(b"01000010010111010100000000000110", b"11000001000100110111100010111000"), -- -64.5295 + 55.3125 = -9.21697
	(b"01000010100001111111111010011110", b"00000000000000000000000000000000"),
	(b"11000010101011011010011011110000", b"11000001100101101010000101001000"), -- 67.9973 + -86.826 = -18.8288
	(b"01000010101100000000000010010000", b"00000000000000000000000000000000"),
	(b"11000010100000100110100011110100", b"01000001101101100101111001110000"), -- 88.0011 + -65.205 = 22.7961
	(b"01000010100011011110000001001111", b"00000000000000000000000000000000"),
	(b"01000000001011010101110110100000", b"01000010100100110100101100111100"), -- 70.9381 + 2.70884 = 73.6469
	(b"01000001010011010100011110111000", b"00000000000000000000000000000000"),
	(b"11000000011101100011010101000000", b"01000001000011111011101001101000"), -- 12.83 + -3.847 = 8.98301
	(b"01000010001010000001000101011011", b"00000000000000000000000000000000"),
	(b"01000010011001010000000111100000", b"01000010110001101000100110011110"), -- 42.0169 + 57.2518 = 99.2688
	(b"11000010101111101001001010011011", b"00000000000000000000000000000000"),
	(b"00111111001100110011010010000000", b"11000010101111010010110000110010"), -- -95.2863 + 0.70002 = -94.5863
	(b"11000010100110011010001110101010", b"00000000000000000000000000000000"),
	(b"11000010100110100010101001100100", b"11000011000110011110011100000111"), -- -76.8197 + -77.0828 = -153.902
	(b"01000001101101010000110111101000", b"00000000000000000000000000000000"),
	(b"11000010001000001011100110111101", b"11000001100011000110010110010010"), -- 22.6318 + -40.1814 = -17.5496
	(b"10111111111111011000000101000000", b"00000000000000000000000000000000"),
	(b"01000000100110110010001011100000", b"01000000001101111000010100100000"), -- -1.98051 + 4.84801 = 2.8675
	(b"11000001001010111101101111011000", b"00000000000000000000000000000000"),
	(b"11000001100011100010000110110100", b"11000001111001000000111110100000"), -- -10.7412 + -17.7665 = -28.5076
	(b"11000000110010011001011101010000", b"00000000000000000000000000000000"),
	(b"01000010100011100110001100111100", b"01000010100000011100100111000111"), -- -6.29972 + 71.1938 = 64.8941
	(b"11000001110110000000111000010000", b"00000000000000000000000000000000"),
	(b"01000010100110011011010001111100", b"01000010010001110110000111110000"), -- -27.0069 + 76.8525 = 49.8456
	(b"01000001101111000111000000110100", b"00000000000000000000000000000000"),
	(b"01000000000101101110011011000000", b"01000001110011110100110100001100"), -- 23.5548 + 2.35783 = 25.9126
	(b"11000001110101000101111111001000", b"00000000000000000000000000000000"),
	(b"11000010000011000111101000100100", b"11000010011101101010101000001000"), -- -26.5468 + -35.1193 = -61.666
	(b"11000001110011111110100101010100", b"00000000000000000000000000000000"),
	(b"01000010100110001110110001110100", b"01000010010010011110010000111110"), -- -25.9889 + 76.4618 = 50.4729
	(b"11000010100001110100000110111010", b"00000000000000000000000000000000"),
	(b"01000010010000101011000110010100", b"11000001100101111010001111000000"), -- -67.6284 + 48.6734 = -18.955
	(b"01000010010100110011001010001110", b"00000000000000000000000000000000"),
	(b"11000010101110010110110011010100", b"11000010000111111010011100011010"), -- 52.7994 + -92.7126 = -39.9132
	(b"01000010100101001011001100011010", b"00000000000000000000000000000000"),
	(b"01000010100111110101101100010000", b"01000011000110100000011100010101"), -- 74.3498 + 79.6779 = 154.028
	(b"01000010001011000111110100101111", b"00000000000000000000000000000000"),
	(b"01000001111001000010000010000000", b"01000010100011110100011010111000"), -- 43.1222 + 28.5159 = 71.6381
	(b"11000010011010000110001011101110", b"00000000000000000000000000000000"),
	(b"01000010011011001011001111110000", b"00111111100010100010000001000000"), -- -58.0966 + 59.1757 = 1.07911
	(b"11000001000101111001111001000000", b"00000000000000000000000000000000"),
	(b"01000010100111000111011000110100", b"01000010100010011000001001101100"), -- -9.47614 + 78.2309 = 68.7547
	(b"11000010100010001011010100100000", b"00000000000000000000000000000000"),
	(b"01000010110000110001000101100000", b"01000001111010010111000100000000"), -- -68.3538 + 97.5339 = 29.1802
	(b"01000010011001010101011100000010", b"00000000000000000000000000000000"),
	(b"11000010100011101010000010101000", b"11000001010111111010100100111000"), -- 57.335 + -71.3138 = -13.9788
	(b"01000010100010100111011000101110", b"00000000000000000000000000000000"),
	(b"01000001011000101100111011100000", b"01000010101001101101000000001010"), -- 69.2308 + 14.1755 = 83.4063
	(b"11000010010101100100011001001110", b"00000000000000000000000000000000"),
	(b"01000001110111001111111110111100", b"11000001110011111000110011100000"), -- -53.5687 + 27.6249 = -25.9438
	(b"01000001000101110101100001110000", b"00000000000000000000000000000000"),
	(b"10111110111100101100100100000000", b"01000001000011111100001000101000"), -- 9.45909 + -0.47419 = 8.9849
	(b"01000010011011100001111100001000", b"00000000000000000000000000000000"),
	(b"10111111100110011010010011000000", b"01000010011010010101000111100010"), -- 59.5303 + -1.20034 = 58.33
	(b"01000001111010100110010110100000", b"00000000000000000000000000000000"),
	(b"11000000101010011001011010110000", b"01000001101111111111111111110100"), -- 29.2996 + -5.29964 = 24
	(b"11000001110111110010010100100000", b"00000000000000000000000000000000"),
	(b"01000010010101100000101110111001", b"01000001110011001111001001010010"), -- -27.8931 + 53.5114 = 25.6183
	(b"11000010001111100011010100000100", b"00000000000000000000000000000000"),
	(b"01000010000000001100000000100000", b"11000001011101011101001110010000"), -- -47.5518 + 32.1876 = -15.3642
	(b"11000010000001110010110001001010", b"00000000000000000000000000000000"),
	(b"01000010101100101000000110111010", b"01000010010111011101011100101010"), -- -33.7933 + 89.2534 = 55.4601
	(b"01000001111000111010000010011000", b"00000000000000000000000000000000"),
	(b"11000010100011100001101101000010", b"11000010001010100110011000111000"), -- 28.4534 + -71.0532 = -42.5998
	(b"11000001100110101100100101101000", b"00000000000000000000000000000000"),
	(b"11000010101000100011111011001110", b"11000010110010001111000100101000"), -- -19.3483 + -81.1227 = -100.471
	(b"11000010101111011111110110000110", b"00000000000000000000000000000000"),
	(b"01000000100010001101011101110000", b"11000010101101010111000000001111"), -- -94.9952 + 4.2763 = -90.7189
	(b"11000010011011101100010111101010", b"00000000000000000000000000000000"),
	(b"11000010101111011000111010001010", b"11000011000110100111100011000000"), -- -59.6933 + -94.7784 = -154.472
	(b"11000010011001101010000111000100", b"00000000000000000000000000000000"),
	(b"01000010011010001100100000011000", b"00111111000010011001010100000000"), -- -57.658 + 58.1954 = 0.53743
	(b"11000001011011101110110111010000", b"00000000000000000000000000000000"),
	(b"11000010010011000100101001000000", b"11000010100001000000001011011010"), -- -14.9331 + -51.0725 = -66.0056
	(b"01000010110000000000010111001111", b"00000000000000000000000000000000"),
	(b"01000010000111100011100011001011", b"01000011000001111001000100011010"), -- 96.0113 + 39.5555 = 135.567
	(b"01000001100110001001000100010100", b"00000000000000000000000000000000"),
	(b"01000010011011001000110001100001", b"01000010100111000110101001110110"), -- 19.0708 + 59.1371 = 78.2079
	(b"11000010011000000000000111011000", b"00000000000000000000000000000000"),
	(b"11000010100100001110010100111000", b"11000011000000000111001100010010"), -- -56.0018 + -72.4477 = -128.449
	(b"11000010101011001000011101101010", b"00000000000000000000000000000000"),
	(b"01000010000111110111010010110000", b"11000010001110011001101000100100"), -- -86.2645 + 39.864 = -46.4005
	(b"01000010000110001001101111010100", b"00000000000000000000000000000000"),
	(b"01000010100110110001100111101110", b"01000010111001110110011111011000"), -- 38.1522 + 77.5506 = 115.703
	(b"11000010010101001000101100111010", b"00000000000000000000000000000000"),
	(b"01000010100010100001110011100001", b"01000001011111101011101000100000"), -- -53.136 + 69.0564 = 15.9204
	(b"01000010101000000010110010000100", b"00000000000000000000000000000000"),
	(b"11000010101101010111110011011010", b"11000001001010101000001010110000"), -- 80.0869 + -90.7439 = -10.6569
	(b"01000010101010100001001100100000", b"00000000000000000000000000000000"),
	(b"11000001011110001100011100111000", b"01000010100010101111101000111001"), -- 85.0374 + -15.5486 = 69.4887
	(b"01000010100100010000000111111010", b"00000000000000000000000000000000"),
	(b"01000010101000001001100000000111", b"01000011000110001100110100000000"), -- 72.5039 + 80.2969 = 152.801
	(b"01000001011100101011110101000000", b"00000000000000000000000000000000"),
	(b"01000010100110010110000101101001", b"01000010101101111011100100010001"), -- 15.1712 + 76.6903 = 91.8615
	(b"11000000010111000011110111000000", b"00000000000000000000000000000000"),
	(b"11000010001110001011011101011000", b"11000010010001100111101100110100"), -- -3.44127 + -46.179 = -49.6203
	(b"01000010101101001000001011101000", b"00000000000000000000000000000000"),
	(b"01000010101111000001000010111101", b"01000011001110000100100111010010"), -- 90.2557 + 94.0327 = 184.288
	(b"01000000100111110011000100000000", b"00000000000000000000000000000000"),
	(b"11000010110000111111011010101110", b"11000010101110100000001110011110"), -- 4.97473 + -97.9818 = -93.0071
	(b"11000010100011001011111011111111", b"00000000000000000000000000000000"),
	(b"01000010010011000111010011110101", b"11000001100110100001001000010010"), -- -70.373 + 51.1142 = -19.2588
	(b"01000010110000000101110110010010", b"00000000000000000000000000000000"),
	(b"01000010000101010101101011010101", b"01000011000001011000010101111110"), -- 96.1828 + 37.3387 = 133.521
	(b"01000001111011010011110110110000", b"00000000000000000000000000000000"),
	(b"11000010001110001101110010110000", b"11000001100001000111101110110000"), -- 29.6551 + -46.2155 = -16.5604
	(b"11000001111100000000101000010100", b"00000000000000000000000000000000"),
	(b"11000010101000000011111001111001", b"11000010110111000100000011111110"), -- -30.0049 + -80.122 = -110.127
	(b"01000001111011100000001111100100", b"00000000000000000000000000000000"),
	(b"01000010001010100111100011010000", b"01000010100100001011110101100001"), -- 29.7519 + 42.618 = 72.3699
	(b"11000010101100111110011000101101", b"00000000000000000000000000000000"),
	(b"11000000000010000011011101000000", b"11000010101110000010011111100111"), -- -89.9496 + -2.12837 = -92.0779
	(b"11000001010101110000001010000000", b"00000000000000000000000000000000"),
	(b"11000010000000000111110111000000", b"11000010001101100011111001100000"), -- -13.4381 + -32.1228 = -45.5609
	(b"11000010101001011110101100010100", b"00000000000000000000000000000000"),
	(b"01000010110001111111010100011100", b"01000001100010000010100000100000"), -- -82.9591 + 99.9787 = 17.0196
	(b"11000000001111011101111110100000", b"00000000000000000000000000000000"),
	(b"01000001001110000000000001000000", b"01000001000010001000100001011000"), -- -2.96677 + 11.5001 = 8.53329
	(b"01000010101110101111010000101010", b"00000000000000000000000000000000"),
	(b"01000010100101000111011100010110", b"01000011001001111011010110100000"), -- 93.4769 + 74.2326 = 167.709
	(b"11000010100000010000100010101110", b"00000000000000000000000000000000"),
	(b"11000010011100111111100101011000", b"11000010111110110000010101011010"), -- -64.517 + -60.9935 = -125.51
	(b"01000010011010001111100001011011", b"00000000000000000000000000000000"),
	(b"01000010010111001100001010100000", b"01000010111000101101110101111110"), -- 58.2425 + 55.1901 = 113.433
	(b"01000010100011100000101010101000", b"00000000000000000000000000000000"),
	(b"01000010001010110000011101000010", b"01000010111000111000111001001001"), -- 71.0208 + 42.7571 = 113.778
	(b"11000010100111001011111110001001", b"00000000000000000000000000000000"),
	(b"01000010101111111101010110011110", b"01000001100011000101100001010100"), -- -78.3741 + 95.9172 = 17.5431
	(b"01000010010100010011110101001100", b"00000000000000000000000000000000"),
	(b"01000010100001011100100011111000", b"01000010111011100110011110011110"), -- 52.3099 + 66.8925 = 119.202
	(b"11000010100100010111100111100000", b"00000000000000000000000000000000"),
	(b"11000001100110000101000011111100", b"11000010101101111000111000011111"), -- -72.738 + -19.0395 = -91.7776
	(b"11000001001011100010011000110000", b"00000000000000000000000000000000"),
	(b"11000010010000100100101010001100", b"11000010011011011101010000011000"), -- -10.8843 + -48.5728 = -59.4571
	(b"11000001101001101100000010110100", b"00000000000000000000000000000000"),
	(b"11000001010000001011001111001000", b"11000010000000111000110101001100"), -- -20.8441 + -12.0439 = -32.888
	(b"11000001111110101101000111110000", b"00000000000000000000000000000000"),
	(b"11000001110101111101010100001000", b"11000010011010010101001101111100"), -- -31.3525 + -26.979 = -58.3315
	(b"11000010011110010000001011010000", b"00000000000000000000000000000000"),
	(b"11000010101010101001100101111101", b"11000011000100111000110101110010"), -- -62.2527 + -85.2998 = -147.553
	(b"01000010011000011001010111101100", b"00000000000000000000000000000000"),
	(b"11000010110000101000110001001101", b"11000010001000111000001010101110"), -- 56.3964 + -97.274 = -40.8776
	(b"01000010100100011110010101010010", b"00000000000000000000000000000000"),
	(b"11000010011000010010110111000001", b"01000001100001010011100111000110"), -- 72.9479 + -56.2947 = 16.6532
	(b"01000010100011101001101100010010", b"00000000000000000000000000000000"),
	(b"00111111100111001011111001000000", b"01000010100100010000111000001011"), -- 71.3029 + 1.22456 = 72.5274
	(b"01000001101100001101010011100100", b"00000000000000000000000000000000"),
	(b"11000010100000010000110101000000", b"11000010001010011011000000001110"), -- 22.104 + -64.5259 = -42.4219
	(b"01000010001011101000000111110101", b"00000000000000000000000000000000"),
	(b"11000000111110011100001010010000", b"01000010000011110100100110100011"), -- 43.6269 + -7.805 = 35.8219
	(b"01000001100010000001010110100000", b"00000000000000000000000000000000"),
	(b"11000010011001011001100001111100", b"11000010001000011000110110101100"), -- 17.0106 + -57.3989 = -40.3884
	(b"11000010100011110110011000011110", b"00000000000000000000000000000000"),
	(b"01000010100100000000110011100100", b"00111110101001101100011000000000"), -- -71.6994 + 72.0252 = 0.325729
	(b"11000010000100011011010000110000", b"00000000000000000000000000000000"),
	(b"01000010100100011010100111000110", b"01000010000100011001111101011100"), -- -36.426 + 72.8316 = 36.4056
	(b"11000001011010011011111100010000", b"00000000000000000000000000000000"),
	(b"11000001010110101000100010011000", b"11000001111000100010001111010100"), -- -14.6091 + -13.6583 = -28.2675
	(b"10111111000000110101010010000000", b"00000000000000000000000000000000"),
	(b"11000010100010011110111101110100", b"11000010100010101111011000011101"), -- -0.513008 + -68.9677 = -69.4807
	(b"11000010100100100001000011110100", b"00000000000000000000000000000000"),
	(b"01000010101110010011010111111100", b"01000001100111001001010000100000"), -- -73.0331 + 92.6054 = 19.5723
	(b"11000001100101110010010000000000", b"00000000000000000000000000000000"),
	(b"11000010000101100110101100011111", b"11000010011000011111110100011111"), -- -18.8926 + -37.6046 = -56.4972
	(b"11000001100011011011100111110100", b"00000000000000000000000000000000"),
	(b"01000010101110111011100111011111", b"01000010100110000100101101100010"), -- -17.7158 + 93.863 = 76.1472
	(b"11000010100111101001011110000101", b"00000000000000000000000000000000"),
	(b"01000010011101101110000001010011", b"11000001100011001001110101101110"), -- -79.2959 + 61.7191 = -17.5769
	(b"11000001100101000111001010010000", b"00000000000000000000000000000000"),
	(b"11000010010001101100111010010100", b"11000010100010001000001111101110"), -- -18.5559 + -49.7017 = -68.2577
	(b"01000010001111001100001110101000", b"00000000000000000000000000000000"),
	(b"11000010100101000111001100010100", b"11000001110110000100010100000000"), -- 47.1911 + -74.2248 = -27.0337
	(b"11000001001001110011000111110000", b"00000000000000000000000000000000"),
	(b"11000010100011011100011111100010", b"11000010101000101010111000100000"), -- -10.4497 + -70.8904 = -81.3401
	(b"01000010010110100110001101001010", b"00000000000000000000000000000000"),
	(b"11000010011111011000001000110100", b"11000001000011000111101110101000"), -- 54.597 + -63.3772 = -8.78019
	(b"11000010101001001110010110001100", b"00000000000000000000000000000000"),
	(b"01000001001110011111110001101000", b"11000010100011011010010111111111"), -- -82.4483 + 11.6241 = -70.8242
	(b"01000010011001011010010010000100", b"00000000000000000000000000000000"),
	(b"01000010101101000010000101000100", b"01000011000100110111100111000011"), -- 57.4107 + 90.065 = 147.476
	(b"00111110111111001011111000000000", b"00000000000000000000000000000000"),
	(b"01000001111010101001000010010000", b"01000001111011101000001110001000"), -- 0.493637 + 29.3206 = 29.8142
	(b"01000010100011100111011111011000", b"00000000000000000000000000000000"),
	(b"01000010001010111110011000101000", b"01000010111001000110101011101100"), -- 71.2341 + 42.9748 = 114.209
	(b"11000010100111101111111100100010", b"00000000000000000000000000000000"),
	(b"01000001111110101111001010000000", b"11000010010000001000010100000100"), -- -79.4983 + 31.3684 = -48.1299
	(b"11000001101101011000101001011100", b"00000000000000000000000000000000"),
	(b"01000010000001110000010010011100", b"01000001001100001111110110111000"), -- -22.6926 + 33.7545 = 11.0619
	(b"01000010000010000101111100101100", b"00000000000000000000000000000000"),
	(b"11000010100000011110000001100110", b"11000001111101101100001101000000"), -- 34.0929 + -64.9383 = -30.8453
	(b"11000010011010111010101010000000", b"00000000000000000000000000000000"),
	(b"11000001111101000110010100011000", b"11000010101100101110111010000110"), -- -58.9165 + -30.5494 = -89.4659
	(b"01000010010101010010011010000100", b"00000000000000000000000000000000"),
	(b"11000010101011110010111100001010", b"11000010000010010011011110010000"), -- 53.2876 + -87.5919 = -34.3043
	(b"11000010000000101001101111000110", b"00000000000000000000000000000000"),
	(b"01000010000110111110111101101100", b"01000000110010101001110100110000"), -- -32.6521 + 38.9838 = 6.33169
	(b"11000010011101110100001011110000", b"00000000000000000000000000000000"),
	(b"01000010110001111110010111010100", b"01000010000110001000100010111000"), -- -61.8154 + 99.9489 = 38.1335
	(b"01000001111111001110011101101000", b"00000000000000000000000000000000"),
	(b"01000001100100001010011111001000", b"01000010010001101100011110011000"), -- 31.613 + 18.0819 = 49.6949
	(b"01000001011110110101010001101000", b"00000000000000000000000000000000"),
	(b"01000010101000000000101101001100", b"01000010101111110111010111011001"), -- 15.7081 + 80.0221 = 95.7302
	(b"01000010100001111000101001000101", b"00000000000000000000000000000000"),
	(b"11000010100101011011111101010110", b"11000000111000110101000100010000"), -- 67.7701 + -74.8737 = -7.10365
	(b"11000010101110001111010100001011", b"00000000000000000000000000000000"),
	(b"11000001010110100000000011001000", b"11000010110101000011010100100100"), -- -92.4786 + -13.6252 = -106.104
	(b"01000010010001111010010010110100", b"00000000000000000000000000000000"),
	(b"11000010011111101000001101011000", b"11000001010110110111101010010000"), -- 49.9108 + -63.6283 = -13.7174
	(b"01000010101110011011000110011010", b"00000000000000000000000000000000"),
	(b"11000010001110111001101000001000", b"01000010001101111100100100101100"), -- 92.8469 + -46.9004 = 45.9465
	(b"11000010101001000010111101000010", b"00000000000000000000000000000000"),
	(b"01000001101101001010000111000000", b"11000010011011100000110110100100"), -- -82.0923 + 22.579 = -59.5133
	(b"01000010100011010101010110001100", b"00000000000000000000000000000000"),
	(b"01000001111110101111111000100100", b"01000010110011000001010100010101"), -- 70.6671 + 31.3741 = 102.041
	(b"01000001010111001100010110010000", b"00000000000000000000000000000000"),
	(b"01000010101101011001111001101000", b"01000010110100010011011100011010"), -- 13.7982 + 90.8094 = 104.608
	(b"11000001100000011001011010110000", b"00000000000000000000000000000000"),
	(b"01000010100100001110010110001101", b"01000010011000001111111111000010"), -- -16.1986 + 72.4483 = 56.2498
	(b"11000010000111110101010001101100", b"00000000000000000000000000000000"),
	(b"01000001001010001011000000100000", b"11000001111010100101000011001000"), -- -39.8324 + 10.543 = -29.2894
	(b"11000010001100110011011101111011", b"00000000000000000000000000000000"),
	(b"00111111110100100000110000000000", b"11000010001011001010011100011011"), -- -44.8042 + 1.64099 = -43.1632
	(b"11000010100010010110111111100010", b"00000000000000000000000000000000"),
	(b"01000010110001010100101000010010", b"01000001111011110110100011000000"), -- -68.7185 + 98.6447 = 29.9261
	(b"11000010000011000011000000001000", b"00000000000000000000000000000000"),
	(b"01000010100111001011111110111100", b"01000010001011010100111101110000"), -- -35.0469 + 78.3745 = 43.3276
	(b"11000001110110001101100001010100", b"00000000000000000000000000000000"),
	(b"01000010001000101011000110101111", b"01000001010110010001011000010100"), -- -27.1056 + 40.6735 = 13.5679
	(b"11000010101000101111000111011110", b"00000000000000000000000000000000"),
	(b"11000010100100010101110100101000", b"11000011000110100010011110000011"), -- -81.4724 + -72.6819 = -154.154
	(b"11000010100100001100110110110100", b"00000000000000000000000000000000"),
	(b"11000000010101110010101011000000", b"11000010100101111000011100001010"), -- -72.4018 + -3.36198 = -75.7637
	(b"11000010010111101111000001101010", b"00000000000000000000000000000000"),
	(b"11000010101010000001010101010110", b"11000011000010111100011011000110"), -- -55.7348 + -84.0417 = -139.776
	(b"01000010100100111100100100001010", b"00000000000000000000000000000000"),
	(b"01000010001111110000111011000100", b"01000010111100110101000001101100"), -- 73.8927 + 47.7644 = 121.657
	(b"11000001010110110111001100001000", b"00000000000000000000000000000000"),
	(b"11000010001010011001011001110000", b"11000010011000000111001100110010"), -- -13.7156 + -42.3969 = -56.1125
	(b"01000010000111001111110010110111", b"00000000000000000000000000000000"),
	(b"11000001000110100001001011100000", b"01000001111011001110111111111110"), -- 39.2468 + -9.62961 = 29.6172
	(b"11000010100110010101100011110100", b"00000000000000000000000000000000"),
	(b"11000000101011101011011000000000", b"11000010101001000100010001010100"), -- -76.6737 + -5.45972 = -82.1335
	(b"01000010101011011011010011001101", b"00000000000000000000000000000000"),
	(b"11000010101001011000010001111010", b"01000000100000110000010100110000"), -- 86.8531 + -82.7587 = 4.09438
	(b"01000000111010110001010011100000", b"00000000000000000000000000000000"),
	(b"11000010011001101111001010111110", b"11000010010010011001000000100010"), -- 7.3463 + -57.7371 = -50.3908
	(b"11000010001100111010011001001100", b"00000000000000000000000000000000"),
	(b"01000010101011100100001000011010", b"01000010001010001101110111101000"), -- -44.9124 + 87.1291 = 42.2167
	(b"11000010001001101001100111000100", b"00000000000000000000000000000000"),
	(b"11000001101000011000000110011100", b"11000010011101110101101010010010"), -- -41.6502 + -20.1883 = -61.8384
	(b"01000010001111111100110101010000", b"00000000000000000000000000000000"),
	(b"11000010000101010011001000011100", b"01000001001010100110110011010000"), -- 47.9505 + -37.2989 = 10.6516
	(b"01000010100100111101110010101010", b"00000000000000000000000000000000"),
	(b"11000010101111010011011010000000", b"11000001101001010110011101011000"), -- 73.931 + -94.6064 = -20.6755
	(b"11000010100111010101011110010100", b"00000000000000000000000000000000"),
	(b"01000001000110101001111110110000", b"11000010100010100000001110011110"), -- -78.6711 + 9.66399 = -69.0071
	(b"01000010100101111100010101010110", b"00000000000000000000000000000000"),
	(b"11000000011010101100001001000000", b"01000010100100000110111101000100"), -- 75.8854 + -3.66811 = 72.2173
	(b"01000010101111011100011110001001", b"00000000000000000000000000000000"),
	(b"11000010010010011100001010011000", b"01000010001100011100110001111010"), -- 94.8897 + -50.44 = 44.4497
	(b"10111111011111110000111100000000", b"00000000000000000000000000000000"),
	(b"01000001101001100110111110111100", b"01000001100111100111011101000100"), -- -0.996323 + 20.8046 = 19.8082
	(b"11000000111111100101000111100000", b"00000000000000000000000000000000"),
	(b"01000001111110100000010010011000", b"01000001101110100111000000100000"), -- -7.94749 + 31.2522 = 23.3047
	(b"01000010010101001010001100111111", b"00000000000000000000000000000000"),
	(b"01000010001111001101111101110101", b"01000010110010001100000101011010"), -- 53.1594 + 47.2182 = 100.378
	(b"01000010100001001011001110010010", b"00000000000000000000000000000000"),
	(b"11000010001000001110111110001011", b"01000001110100001110111100110010"), -- 66.3507 + -40.2339 = 26.1168
	(b"11000010011011111010110011100101", b"00000000000000000000000000000000"),
	(b"01000010000001111100110010001100", b"11000001110011111100000010110010"), -- -59.9188 + 33.9498 = -25.9691
	(b"11000010010010000010100100001101", b"00000000000000000000000000000000"),
	(b"01000010110000101000011011010100", b"01000010001111001110010010011011"), -- -50.0401 + 97.2633 = 47.2232
	(b"11000010101011100100000111011000", b"00000000000000000000000000000000"),
	(b"01000010110001110101000001100010", b"01000001010010000111010001010000"), -- -87.1286 + 99.657 = 12.5284
	(b"11000010101111010010000110011000", b"00000000000000000000000000000000"),
	(b"01000000101111100010001000000000", b"11000010101100010011111101111000"), -- -94.5656 + 5.94165 = -88.624
	(b"01000010001111110011011011000000", b"00000000000000000000000000000000"),
	(b"01000010101000101001011010010100", b"01000011000000010001100011111010"), -- 47.8035 + 81.2941 = 129.098
	(b"11000010101111000101110101010010", b"00000000000000000000000000000000"),
	(b"01000001110111111110100101010000", b"11000010100001000110001011111110"), -- -94.1823 + 27.9889 = -66.1933
	(b"11000010101100101110100111110000", b"00000000000000000000000000000000"),
	(b"11000010010100101010001101010000", b"11000011000011100001110111001100"), -- -89.4569 + -52.6595 = -142.116
	(b"01000010100100111110000111111000", b"00000000000000000000000000000000"),
	(b"11000010001110111110101110101100", b"01000001110101111011000010001000"), -- 73.9413 + -46.9801 = 26.9612
	(b"11000010101100000101011100001100", b"00000000000000000000000000000000"),
	(b"01000001100010011001010010010000", b"11000010100011011111000111101000"), -- -88.17 + 17.1975 = -70.9725
	(b"11000010100010101110111001001000", b"00000000000000000000000000000000"),
	(b"01000010010111101011001100001010", b"11000001010111001010011000011000"), -- -69.4654 + 55.6748 = -13.7906
	(b"01000001100111001011000100011000", b"00000000000000000000000000000000"),
	(b"01000010001011100010111001011000", b"01000010011111001000011011100100"), -- 19.5865 + 43.5453 = 63.1317
	(b"01000010100001011001000101010010", b"00000000000000000000000000000000"),
	(b"01000010011110010010011010011100", b"01000011000000010001001001010000"), -- 66.7838 + 62.2877 = 129.072
	(b"00111111010100010111010010000000", b"00000000000000000000000000000000"),
	(b"11000010010010011010010000101100", b"11000010010001100101111001011010"), -- 0.818184 + -50.4103 = -49.5921
	(b"01000001100001110001011010000100", b"00000000000000000000000000000000"),
	(b"01000010101101100101001000101110", b"01000010110110000001011111001111"), -- 16.886 + 91.1605 = 108.047
	(b"01000010010101001000100100000100", b"00000000000000000000000000000000"),
	(b"01000001110100001111101111101000", b"01000010100111101000001101111100"), -- 53.1338 + 26.123 = 79.2568
	(b"11000010101001101110000000010001", b"00000000000000000000000000000000"),
	(b"11000010101000101010001000101110", b"11000011001001001100000100100000"), -- -83.4376 + -81.3168 = -164.754
	(b"01000010100000011110100110011110", b"00000000000000000000000000000000"),
	(b"11000001011000100001110001101000", b"01000010010010110100110000100010"), -- 64.9563 + -14.1319 = 50.8243
	(b"11000010100111000011000000101010", b"00000000000000000000000000000000"),
	(b"11000010110000001111111101010111", b"11000011001011101001011111000000"), -- -78.0941 + -96.4987 = -174.593
	(b"01000000101010010100011010000000", b"00000000000000000000000000000000"),
	(b"01000010010101100011000100011111", b"01000010011010110101100111101111"), -- 5.28986 + 53.548 = 58.8378
	(b"01000010101011010100111010011100", b"00000000000000000000000000000000"),
	(b"11000000110001101000111001000000", b"01000010101000001110010110111000"), -- 86.6535 + -6.20486 = 80.4487
	(b"01000010010100111100011011101100", b"00000000000000000000000000000000"),
	(b"01000010101101001101111101110011", b"01000011000011110110000101110100"), -- 52.9443 + 90.4364 = 143.381
	(b"01000010010011011100010111010000", b"00000000000000000000000000000000"),
	(b"11000010001000111111011110110100", b"01000001001001110011100001110000"), -- 51.4432 + -40.9919 = 10.4513
	(b"11000010101101100111010110001000", b"00000000000000000000000000000000"),
	(b"11000010001101010000001001011100", b"11000011000010000111101101011011"), -- -91.2296 + -45.2523 = -136.482
	(b"11000000101011001100111001100000", b"00000000000000000000000000000000"),
	(b"01000010100101001110100100010101", b"01000010100010100001110000101111"), -- -5.40019 + 74.4552 = 69.055
	(b"11000010011111101100010111001100", b"00000000000000000000000000000000"),
	(b"01000001111110011110110001110000", b"11000010000000011100111110010100"), -- -63.6932 + 31.2404 = -32.4527
	(b"11000010100001100111111111100000", b"00000000000000000000000000000000"),
	(b"01000010101111111111100100001101", b"01000001111001011110010010110100"), -- -67.2498 + 95.9864 = 28.7367
	(b"11000010001010101001011111110011", b"00000000000000000000000000000000"),
	(b"01000001011100110011011000000000", b"11000001110110111001010011100110"), -- -42.6484 + 15.2007 = -27.4477
	(b"01000010010001011010000000101010", b"00000000000000000000000000000000"),
	(b"01000010100010111110100011010110", b"01000010111011101011100011101011"), -- 49.4064 + 69.9548 = 119.361
	(b"01000001111011000110110100010000", b"00000000000000000000000000000000"),
	(b"00111111111111010011011001000000", b"01000001111111000100000001110100"), -- 29.5533 + 1.97822 = 31.5315
	(b"01000010100101010001110111010001", b"00000000000000000000000000000000"),
	(b"01000001000000100010011001101000", b"01000010101001010110001010011110"), -- 74.5582 + 8.13438 = 82.6926
	(b"10111111011100011011000000000000", b"00000000000000000000000000000000"),
	(b"11000010110000000110010100110111", b"11000010110000100100100010010111"), -- -0.944092 + -96.1977 = -97.1418
	(b"01000010000110100010101100011001", b"00000000000000000000000000000000"),
	(b"11000010101010110101011010010101", b"11000010001111001000001000010001"), -- 38.5421 + -85.6691 = -47.127
	(b"01000001111010001001001111101000", b"00000000000000000000000000000000"),
	(b"01000001000000010011101111001000", b"01000010000101001001100011100110"), -- 29.0722 + 8.0771 = 37.1493
	(b"11000010110001100100001000100100", b"00000000000000000000000000000000"),
	(b"01000010100001100000111010001000", b"11000010000000000110011100111000"), -- -99.1292 + 67.0284 = -32.1008
	(b"11000001110111100111011100001000", b"00000000000000000000000000000000"),
	(b"11000010000101011010101011110100", b"11000010100000100111001100111100"), -- -27.8081 + -37.4169 = -65.2251
	(b"01000010100011000001101110001010", b"00000000000000000000000000000000"),
	(b"01000010100010001000011001100000", b"01000011000010100101000011110101"), -- 70.0538 + 68.2625 = 138.316
	(b"01000010010101110110011101000111", b"00000000000000000000000000000000"),
	(b"11000010000111010100010110101100", b"01000001011010001000011001101100"), -- 53.8509 + -39.318 = 14.5328
	(b"11000010101100001111111111101100", b"00000000000000000000000000000000"),
	(b"11000001100010001011011100110100", b"11000010110100110010110110111001"), -- -88.4998 + -17.0895 = -105.589
	(b"11000010100011111010110100101000", b"00000000000000000000000000000000"),
	(b"11000001101011010000111110011100", b"11000010101110101111000100001111"), -- -71.8382 + -21.6326 = -93.4708
	(b"01000010100110100000001100100100", b"00000000000000000000000000000000"),
	(b"01000001011000011010010100000000", b"01000010101101100011011111000100"), -- 77.0061 + 14.1028 = 91.1089
	(b"01000010101111110111100011101010", b"00000000000000000000000000000000"),
	(b"11000001001100111011110111011000", b"01000010101010010000000100101111"), -- 95.7362 + -11.2338 = 84.5023
	(b"11000010100001011001011110101110", b"00000000000000000000000000000000"),
	(b"01000001000101110101001010110000", b"11000010011001010101101010110000"), -- -66.7962 + 9.45769 = -57.3386
	(b"01000010011111100100110110000100", b"00000000000000000000000000000000"),
	(b"01000010001000110011101011000100", b"01000010110100001100010000100100"), -- 63.5757 + 40.8074 = 104.383
	(b"11000010100100100101000001001110", b"00000000000000000000000000000000"),
	(b"01000010100111000011100101001110", b"01000000100111101001000000000000"), -- -73.1568 + 78.1119 = 4.95508
	(b"01000010100011001110101101110110", b"00000000000000000000000000000000"),
	(b"11000001000110010100111100001000", b"01000010011100111000001100101010"), -- 70.4599 + -9.58179 = 60.8781
	(b"01000001100110100010111011000100", b"00000000000000000000000000000000"),
	(b"11000010011100101001000010000100", b"11000010001001010111100100100010"), -- 19.2728 + -60.6411 = -41.3683
	(b"01000010101111011010000001010010", b"00000000000000000000000000000000"),
	(b"11000010101000000111011110010100", b"01000001011010010100010111110000"), -- 94.8131 + -80.2336 = 14.5796
	(b"11000010001011000011010111111100", b"00000000000000000000000000000000"),
	(b"11000000101101000010000011100000", b"11000010010000101011101000011000"), -- -43.0527 + -5.62901 = -48.6817
	(b"01000001001111110101101010111000", b"00000000000000000000000000000000"),
	(b"11000010001000110101100111101100", b"11000001111001110000011001111100"), -- 11.9596 + -40.8378 = -28.8782
	(b"11000010001110111111101101011100", b"00000000000000000000000000000000"),
	(b"01000010000001110010100100011010", b"11000001010100110100100100001000"), -- -46.9955 + 33.7901 = -13.2053
	(b"01000001100011010001011110100000", b"00000000000000000000000000000000"),
	(b"01000010010010100100001001011100", b"01000010100010000110011100010110"), -- 17.6365 + 50.5648 = 68.2013
	(b"11000010011101101100011111101100", b"00000000000000000000000000000000"),
	(b"11000010100101001011001100100100", b"11000011000010000000101110001101"), -- -61.6952 + -74.3499 = -136.045
	(b"01000010101101111111011100110100", b"00000000000000000000000000000000"),
	(b"11000010011111010010110011010010", b"01000001111001011000001100101100"), -- 91.9828 + -63.2938 = 28.689
	(b"10111110111000110111101000000000", b"00000000000000000000000000000000"),
	(b"11000010100001000100001001001110", b"11000010100001010010010111001000"), -- -0.44429 + -66.1295 = -66.5738
	(b"11000010110001100111111000001100", b"00000000000000000000000000000000"),
	(b"01000010010100000000011100001111", b"11000010001111001111010100001001"), -- -99.2462 + 52.0069 = -47.2393
	(b"01000010000010101111001000000000", b"00000000000000000000000000000000"),
	(b"11000010000011001011000000010010", b"10111110110111110000100100000000"), -- 34.7363 + -35.1719 = -0.435616
	(b"01000000111111101000111010000000", b"00000000000000000000000000000000"),
	(b"11000010101111000110110010011000", b"11000010101011001000001110110000"), -- 7.9549 + -94.2121 = -86.2572
	(b"11000001010101101110010111111000", b"00000000000000000000000000000000"),
	(b"11000010101010111001001010000100", b"11000010110001100110111101000011"), -- -13.4311 + -85.7862 = -99.2173
	(b"01000010100010000000101110010010", b"00000000000000000000000000000000"),
	(b"11000010101001011000001001101000", b"11000001011010111011011010110000"), -- 68.0226 + -82.7547 = -14.7321
	(b"01000010011000110011010010000100", b"00000000000000000000000000000000"),
	(b"01000001100011010000111001011000", b"01000010100101001101110111011000"), -- 56.8013 + 17.632 = 74.4333
	(b"01000010110001101110111001001110", b"00000000000000000000000000000000"),
	(b"11000001110101000111111100011000", b"01000010100100011100111010001000"), -- 99.4654 + -26.5621 = 72.9034
	(b"01000010101100111111101000101001", b"00000000000000000000000000000000"),
	(b"11000010100110001100001001110000", b"01000001010110011011110111001000"), -- 89.9886 + -76.3798 = 13.6088
	(b"01000010010101101000111000100001", b"00000000000000000000000000000000"),
	(b"11000001000110110110000001101000", b"01000010001011111011011000000111"), -- 53.6388 + -9.71104 = 43.9278
	(b"11000010010011010010111000000100", b"00000000000000000000000000000000"),
	(b"11000000000101110010000101000000", b"11000010010101101010000000011000"), -- -51.2949 + -2.3614 = -53.6563
	(b"01000010011011000101100000010100", b"00000000000000000000000000000000"),
	(b"11000010100010000000100111010011", b"11000001000011101110111001001000"), -- 59.086 + -68.0192 = -8.93317
	(b"11000001111010110110011101101000", b"00000000000000000000000000000000"),
	(b"11000010001111001001010001111100", b"11000010100110010010010000011000"), -- -29.4255 + -47.145 = -76.5705
	(b"11000010101111000001000000011010", b"00000000000000000000000000000000"),
	(b"01000010000011001111111001101100", b"11000010011010110010000111001000"), -- -94.0314 + 35.2485 = -58.783
	(b"01000001001111111110110011001000", b"00000000000000000000000000000000"),
	(b"01000001111011111000111011010000", b"01000010001001111100001010011010"), -- 11.9953 + 29.9447 = 41.94
	(b"11000010011111000010101010101110", b"00000000000000000000000000000000"),
	(b"11000010010011110000110001000101", b"11000010111001011001101101111010"), -- -63.0417 + -51.762 = -114.804
	(b"11000000101111011110010010100000", b"00000000000000000000000000000000"),
	(b"01000010011000110101011110111011", b"01000010010010111001101100100111"), -- -5.93416 + 56.8357 = 50.9015
	(b"01000001100111110101101001110100", b"00000000000000000000000000000000"),
	(b"01000010010101100100101110000110", b"01000010100100101111110001100000"), -- 19.9192 + 53.5738 = 73.4929
	(b"01000010001011101010000001100000", b"00000000000000000000000000000000"),
	(b"01000000110000010101011000010000", b"01000010010001101100101100100010"), -- 43.6566 + 6.04176 = 49.6984
	(b"01000000110101001100100000110000", b"00000000000000000000000000000000"),
	(b"01000001100101100000101010101100", b"01000001110010110011110010111000"), -- 6.64944 + 18.7552 = 25.4046
	(b"01000010110000001111000100110010", b"00000000000000000000000000000000"),
	(b"01000010101010101000101000100000", b"01000011001101011011110110101001"), -- 96.4711 + 85.2698 = 181.741
	(b"01000010011001111111101000000100", b"00000000000000000000000000000000"),
	(b"01000010100011101110000110101100", b"01000011000000010110111101010111"), -- 57.9942 + 71.4408 = 129.435
	(b"11000010000100100101001001100100", b"00000000000000000000000000000000"),
	(b"11000010001001000111010010010100", b"11000010100110110110001101111100"), -- -36.5805 + -41.1138 = -77.6943
	(b"01000010011100101000001101000000", b"00000000000000000000000000000000"),
	(b"11000010010000000110101001111100", b"01000001010010000110001100010000"), -- 60.6282 + -48.104 = 12.5242
	(b"11000010100100101100111010101100", b"00000000000000000000000000000000"),
	(b"01000010010110010111111111100000", b"11000001100110000011101011110000"), -- -73.4037 + 54.3749 = -19.0288
	(b"01000001101011100011000010101100", b"00000000000000000000000000000000"),
	(b"01000010101110111100011101110000", b"01000010111001110101001110011011"), -- 21.7738 + 93.8895 = 115.663
	(b"11000010000000011110010111001110", b"00000000000000000000000000000000"),
	(b"11000010010101001000100001111000", b"11000010101010110011011100100011"), -- -32.4744 + -53.1333 = -85.6077
	(b"11000010100111001001100101110100", b"00000000000000000000000000000000"),
	(b"11000010001011111101100110111000", b"11000010111101001000011001010000"), -- -78.2997 + -43.9626 = -122.262
	(b"11000010101001001100101010101010", b"00000000000000000000000000000000"),
	(b"11000001001111000010000110010000", b"11000010101111000100111011011100"), -- -82.3958 + -11.7582 = -94.154
	(b"01000010101100010111001011011000", b"00000000000000000000000000000000"),
	(b"11000010000111001101010110100100", b"01000010010001100001000000001100"), -- 88.7243 + -39.2086 = 49.5157
	(b"01000010001111001010111000101000", b"00000000000000000000000000000000"),
	(b"01000010101110110000101100101101", b"01000011000011001011000100100000"), -- 47.1701 + 93.5218 = 140.692
	(b"11000000100110001111000101010000", b"00000000000000000000000000000000"),
	(b"11000001111010000001100111011000", b"11000010000001110010101100010110"), -- -4.77946 + -29.0126 = -33.7921
	(b"01000010001110011001001010101000", b"00000000000000000000000000000000"),
	(b"01000001110101101110110000010000", b"01000010100100101000010001011000"), -- 46.3932 + 26.8653 = 73.2585
	(b"01000010110001100010100101100101", b"00000000000000000000000000000000"),
	(b"11000000100110011100111001010000", b"01000010101111001000110010000000"), -- 99.0808 + -4.80643 = 94.2744
	(b"11000010100110101110111011101110", b"00000000000000000000000000000000"),
	(b"11000010100011101011011111111010", b"11000011000101001101001101110100"), -- -77.4667 + -71.3593 = -148.826
	(b"01000010101001010011011101110110", b"00000000000000000000000000000000"),
	(b"11000010010011101000101000100100", b"01000001111101111100100110010000"), -- 82.6083 + -51.6349 = 30.9734
	(b"11000010110000010011101101000100", b"00000000000000000000000000000000"),
	(b"10111111110100010100000101000000", b"11000010110001001000000001001001"), -- -96.6158 + -1.6348 = -98.2506
	(b"01000010010111010100100101010000", b"00000000000000000000000000000000"),
	(b"01000010110000101000111111011100", b"01000011000110001001101001000010"), -- 55.3216 + 97.281 = 152.603
	(b"01000010011010010101001010100000", b"00000000000000000000000000000000"),
	(b"01000001001100010101110110111000", b"01000010100010101101010100000111"), -- 58.3307 + 11.0854 = 69.4161
	(b"11000010001111011110011011101000", b"00000000000000000000000000000000"),
	(b"01000010110000011111111010111110", b"01000010010001100001011010010100"), -- -47.4755 + 96.9975 = 49.522
	(b"01000001110100101000011010001000", b"00000000000000000000000000000000"),
	(b"11000010101100110011100010011100", b"11000010011111010010110111110100"), -- 26.3157 + -89.6106 = -63.2949
	(b"01000001101010000110101010010100", b"00000000000000000000000000000000"),
	(b"11000010101001110010010000101000", b"11000010011110100001001100000110"), -- 21.052 + -83.5706 = -62.5186
	(b"11000001100100100101110111110100", b"00000000000000000000000000000000"),
	(b"01000010000111010000000010101111", b"01000001101001111010001101101010"), -- -18.2959 + 39.2507 = 20.9548
	(b"11000010101001101010111100100110", b"00000000000000000000000000000000"),
	(b"11000010001000000010011011111010", b"11000010111101101100001010100011"), -- -83.3421 + -40.0381 = -123.38
	(b"11000010000011000111011110010000", b"00000000000000000000000000000000"),
	(b"11000001000110010001100101000000", b"11000010001100101011110111100000"), -- -35.1168 + -9.56866 = -44.6854
	(b"01000010101011101101001000001110", b"00000000000000000000000000000000"),
	(b"11000010000100101010000000111100", b"01000010010010110000001111100000"), -- 87.4103 + -36.6565 = 50.7538
	(b"01000010100000110001010111000100", b"00000000000000000000000000000000"),
	(b"01000010001111010100101011011100", b"01000010111000011011101100110010"), -- 65.5425 + 47.3231 = 112.866
	(b"01000010100000100100101011111100", b"00000000000000000000000000000000"),
	(b"01000010011111011101010110001100", b"01000011000000001001101011100001"), -- 65.1465 + 63.4585 = 128.605
	(b"11000010100011000100001001001110", b"00000000000000000000000000000000"),
	(b"11000001001110011111110100100000", b"11000010101000111000000111110010"), -- -70.1295 + -11.6243 = -81.7538
	(b"01000010010000000010100010111011", b"00000000000000000000000000000000"),
	(b"01000010011100010011000101010101", b"01000010110110001010110100001000"), -- 48.0398 + 60.2982 = 108.338
	(b"01000010000011001110100100001110", b"00000000000000000000000000000000"),
	(b"11000001000010101000101110001000", b"01000001110101001000110001011000"), -- 35.2276 + -8.65907 = 26.5685
	(b"01000010101101000100000010101101", b"00000000000000000000000000000000"),
	(b"11000001100010101001100010000000", b"01000010100100011001101010001101"), -- 90.1263 + -17.3245 = 72.8019
	(b"11000010100010001101100100010000", b"00000000000000000000000000000000"),
	(b"01000010100011011100011001111110", b"01000000000111011010110111000000"), -- -68.424 + 70.8877 = 2.46373
	(b"11000010000000110000010110011000", b"00000000000000000000000000000000"),
	(b"11000001101010001000111001011000", b"11000010010101110100110011000100"), -- -32.7555 + -21.0695 = -53.825
	(b"01000001001110110000010111001000", b"00000000000000000000000000000000"),
	(b"11000001111000101001110111000000", b"11000001100001010001101011011100"), -- 11.6889 + -28.327 = -16.6381
	(b"11000001000100011100100011001000", b"00000000000000000000000000000000"),
	(b"01000010000011001111111010000100", b"01000001110100010001100010100100"), -- -9.11152 + 35.2486 = 26.137
	(b"11000000000011110110100100100000", b"00000000000000000000000000000000"),
	(b"11000001101001101111011111110100", b"11000001101110001110010100011000"), -- -2.24079 + -20.8711 = -23.1119
	(b"01000001100010101110100011110000", b"00000000000000000000000000000000"),
	(b"11000001100011001100011101000000", b"10111110011011110010100000000000"), -- 17.3637 + -17.5973 = -0.233551
	(b"01000010110000101011110100110000", b"00000000000000000000000000000000"),
	(b"11000010010000011110000000010000", b"01000010010000111001101001010000"), -- 97.3695 + -48.4688 = 48.9007
	(b"01000001011010001000011011010000", b"00000000000000000000000000000000"),
	(b"01000010100010101111010001110010", b"01000010101010000000010101001100"), -- 14.5329 + 69.4774 = 84.0103
	(b"11000010110001101110011110011100", b"00000000000000000000000000000000"),
	(b"11000010001000100011000001000101", b"11000011000010111111111111011111"), -- -99.4524 + -40.5471 = -139.999
	(b"11000010010000010010101010010100", b"00000000000000000000000000000000"),
	(b"11000010100110100000000001001100", b"11000010111110101001010110010110"), -- -48.2916 + -77.0006 = -125.292
	(b"01000010000111101001001010101100", b"00000000000000000000000000000000"),
	(b"01000010000001010110001110000100", b"01000010100100011111101100011000"), -- 39.6432 + 33.3472 = 72.9904
	(b"11000010100111010111101101011110", b"00000000000000000000000000000000"),
	(b"11000001111001010010001000000100", b"11000010110101101100001111011111"), -- -78.741 + -28.6416 = -107.383
	(b"11000001010100011000000111110000", b"00000000000000000000000000000000"),
	(b"01000001000101111100110100001000", b"11000000011001101101001110100000"), -- -13.0942 + 9.48756 = -3.60667
	(b"11000010101101011111101010101110", b"00000000000000000000000000000000"),
	(b"11000010101010000100101101000011", b"11000011001011110010001011111000"), -- -90.9896 + -84.147 = -175.137
	(b"11000010011111001010010011111111", b"00000000000000000000000000000000"),
	(b"01000001110101101001101011100000", b"11000010000100010101011110001111"), -- -63.1611 + 26.8256 = -36.3355
	(b"01000001110011101100101100011000", b"00000000000000000000000000000000"),
	(b"01000010100100011010111001010010", b"01000010110001010110000100011000"), -- 25.8492 + 72.8405 = 98.6896
	(b"01000010101010111001110010010010", b"00000000000000000000000000000000"),
	(b"01000001101101011011110001011000", b"01000010110110010000101110101000"), -- 85.8058 + 22.717 = 108.523
	(b"01000010010100011101010111100000", b"00000000000000000000000000000000"),
	(b"11000010000101010100101010101100", b"01000001011100100010110011010000"), -- 52.4589 + -37.3229 = 15.1359
	(b"11000010101001110011101011111011", b"00000000000000000000000000000000"),
	(b"01000010001101111100010100011000", b"11000010000101101011000011011110"), -- -83.6152 + 45.9425 = -37.6727
	(b"11000010101101110011010110110100", b"00000000000000000000000000000000"),
	(b"01000000111011010001111001000000", b"11000010101010000110001111010000"), -- -91.6049 + 7.40994 = -84.1949
	(b"01000001010000110110100000101000", b"00000000000000000000000000000000"),
	(b"11000001100001110110001101001100", b"11000000100101101011110011100000"), -- 12.2129 + -16.9235 = -4.71056
	(b"11000001111110101010001010100100", b"00000000000000000000000000000000"),
	(b"01000010100101000001100010011100", b"01000010001010101101111111100110"), -- -31.3294 + 74.0481 = 42.7187
	(b"11000010011110001001101101110100", b"00000000000000000000000000000000"),
	(b"01000001100000000111011010000000", b"11000010001110000110000000110100"), -- -62.1518 + 16.0579 = -46.0939
	(b"01000001111010100100000010101000", b"00000000000000000000000000000000"),
	(b"11000010011011001001100001011000", b"11000001111011101111000000001000"), -- 29.2816 + -59.1488 = -29.8672
	(b"01000010110001101000000010010010", b"00000000000000000000000000000000"),
	(b"11000010001011010000001000101000", b"01000010010111111111111011111100"), -- 99.2511 + -43.2521 = 55.999
	(b"01000010001001010011110010111111", b"00000000000000000000000000000000"),
	(b"01000001110001011100111001101000", b"01000010100001000001000111111010"), -- 41.3093 + 24.7258 = 66.0351
	(b"01000010010100100111101010101100", b"00000000000000000000000000000000"),
	(b"11000001100001000010101101101100", b"01000010000100000110010011110110"), -- 52.6198 + -16.5212 = 36.0986
	(b"01000010000000111101110101110110", b"00000000000000000000000000000000"),
	(b"01000010101111001101001111101001", b"01000010111111101100001010100100"), -- 32.9663 + 94.4139 = 127.38
	(b"11000010001000110111101010011000", b"00000000000000000000000000000000"),
	(b"01000010000111110101011010101000", b"10111111100001000111111000000000"), -- -40.8697 + 39.8346 = -1.0351
	(b"01000010110000111010100110011100", b"00000000000000000000000000000000"),
	(b"01000010000101011001100111000100", b"01000011000001110011101100111111"), -- 97.8313 + 37.4002 = 135.231
	(b"11000010011111101101000100000111", b"00000000000000000000000000000000"),
	(b"01000001011101010110000100101000", b"11000010010000010111100010111101"), -- -63.7041 + 15.3362 = -48.3679
	(b"11000010011001100011111110010000", b"00000000000000000000000000000000"),
	(b"01000010100011000010101001100010", b"01000001010010000101010011010000"), -- -57.5621 + 70.0828 = 12.5207
	(b"01000010101011110111010001100100", b"00000000000000000000000000000000"),
	(b"11000000001011011011011001000000", b"01000010101010100000011010110010"), -- 87.7273 + -2.71425 = 85.0131
	(b"11000010011011011011011001011000", b"00000000000000000000000000000000"),
	(b"11000010101101111001001100000110", b"11000011000101110011011100011001"), -- -59.4281 + -91.7872 = -151.215
	(b"01000010100000100001100111001110", b"00000000000000000000000000000000"),
	(b"01000010001010100011011010101000", b"01000010110101110011010100100010"), -- 65.0504 + 42.5534 = 107.604
	(b"11000001111001101110101100000000", b"00000000000000000000000000000000"),
	(b"11000010000000010101010100110000", b"11000010011101001100101010110000"), -- -28.8647 + -32.3332 = -61.1979
	(b"11000010010011110000011010010000", b"00000000000000000000000000000000"),
	(b"01000010100011000111010110000100", b"01000001100100111100100011110000"), -- -51.7564 + 70.2295 = 18.4731
	(b"11000010101110001000111111100100", b"00000000000000000000000000000000"),
	(b"01000010101110110101000000101100", b"00111111101100000001001000000000"), -- -92.281 + 93.6566 = 1.37555
	(b"01000010100111110000100000011101", b"00000000000000000000000000000000"),
	(b"01000010101011101000100011010000", b"01000011001001101100100001110110"), -- 79.5158 + 87.2672 = 166.783
	(b"11000010101000011101100111010110", b"00000000000000000000000000000000"),
	(b"01000000010100111111000011000000", b"11000010100110110011101001010000"), -- -80.9255 + 3.31157 = -77.6139
	(b"11000000001010110010111111100000", b"00000000000000000000000000000000"),
	(b"11000010011011111001011111000000", b"11000010011110100100101010111110"), -- -2.6748 + -59.8982 = -62.573
	(b"11000001001001110100010110001000", b"00000000000000000000000000000000"),
	(b"11000001011010010100101010000000", b"11000001110010000100100000000100"), -- -10.4545 + -14.5807 = -25.0352
	(b"01000010101001110000100100111110", b"00000000000000000000000000000000"),
	(b"01000010010001000001000101110111", b"01000011000001001000100011111101"), -- 83.5181 + 49.0171 = 132.535
	(b"11000010010100100010001100101100", b"00000000000000000000000000000000"),
	(b"11000010100010101100001010110110", b"11000010111100111101010001001100"), -- -52.5343 + -69.3803 = -121.915
	(b"01000010101101000000111101001100", b"00000000000000000000000000000000"),
	(b"01000010110001011110100100000001", b"01000011001111001111110000100110"), -- 90.0299 + 98.9551 = 188.985
	(b"01000001101001101110111011011000", b"00000000000000000000000000000000"),
	(b"11000001110101000100000111001100", b"11000000101101010100101111010000"), -- 20.8666 + -26.5321 = -5.6655
	(b"11000010010000110101100110110000", b"00000000000000000000000000000000"),
	(b"11000010101011000010001110000101", b"11000011000001101110100000101110"), -- -48.8376 + -86.0694 = -134.907
	(b"11000001111100111011101000101000", b"00000000000000000000000000000000"),
	(b"11000001111100001011010101100000", b"11000010011100100011011111000100"), -- -30.4659 + -30.0886 = -60.5545
	(b"11000010100010011110100110011100", b"00000000000000000000000000000000"),
	(b"01000001111011010100010100011000", b"11000010000111010011000010101100"), -- -68.9563 + 29.6587 = -39.2975
	(b"11000001100110010101010100001000", b"00000000000000000000000000000000"),
	(b"01000010101110010001100000011010", b"01000010100100101100001011011000"), -- -19.1665 + 92.5471 = 73.3806
	(b"11000010101001100100111110001100", b"00000000000000000000000000000000"),
	(b"11000010000010110111100001100000", b"11000010111011000000101110111100"), -- -83.1554 + -34.8676 = -118.023
	(b"01000001111001111101110011100000", b"00000000000000000000000000000000"),
	(b"01000010100111111001110101010010", b"01000010110110011001010010001010"), -- 28.9828 + 79.8073 = 108.79
	(b"11000010100000110100101000100100", b"00000000000000000000000000000000"),
	(b"01000010110000001110100111010001", b"01000001111101100111111010110100"), -- -65.6448 + 96.4567 = 30.8119
	(b"11000010100000000011110100101000", b"00000000000000000000000000000000"),
	(b"01000010010010100110010001011000", b"11000001010110000101011111100000"), -- -64.1194 + 50.598 = -13.5215
	(b"11000001001011100000001110011000", b"00000000000000000000000000000000"),
	(b"11000001101110001010110000101000", b"11000010000001111101011011111010"), -- -10.8759 + -23.0841 = -33.9599
	(b"11000010101111100100000010000100", b"00000000000000000000000000000000"),
	(b"01000010100100110100001001100000", b"11000001101010111111100010010000"), -- -95.126 + 73.6296 = -21.4964
	(b"11000010001101101001010101011000", b"00000000000000000000000000000000"),
	(b"11000001000000010101011001000000", b"11000010010101101110101011101000"), -- -45.6458 + -8.08356 = -53.7294
	(b"11000010100100110001001000100000", b"00000000000000000000000000000000"),
	(b"01000001110000010111001010110000", b"11000010010001010110101011101000"), -- -73.5354 + 24.181 = -49.3544
	(b"01000001100101000010100010111100", b"00000000000000000000000000000000"),
	(b"01000010100100000110111111001001", b"01000010101101010111100111111000"), -- 18.5199 + 72.2183 = 90.7382
	(b"01000010101101001000111110010010", b"00000000000000000000000000000000"),
	(b"01000010010111011001110011100100", b"01000011000100011010111100000010"), -- 90.2804 + 55.4032 = 145.684
	(b"01000010011111100101111111110001", b"00000000000000000000000000000000"),
	(b"11000010001110100001000001110100", b"01000001100010001001111011111010"), -- 63.5937 + -46.5161 = 17.0776
	(b"01000010110001001000111001011000", b"00000000000000000000000000000000"),
	(b"01000010000100011101110111110000", b"01000011000001101011111010101000"), -- 98.278 + 36.4667 = 134.745
	(b"11000010001100010101100101000000", b"00000000000000000000000000000000"),
	(b"01000010100101100101001110011110", b"01000001111101101001101111111000"), -- -44.3372 + 75.1633 = 30.8262
	(b"01000001000010011010010101001000", b"00000000000000000000000000000000"),
	(b"01000001110011001011101110010100", b"01000010000010001100011100011100"), -- 8.60285 + 25.5916 = 34.1944
	(b"11000010001011100010100111011100", b"00000000000000000000000000000000"),
	(b"11000010000010000100101000101000", b"11000010100110110011101000000010"), -- -43.5409 + -34.0724 = -77.6133
	(b"11000010011110111101000101010101", b"00000000000000000000000000000000"),
	(b"01000010011111110101101011001100", b"00111111011000100101110111000000"), -- -62.9544 + 63.8387 = 0.884243
	(b"01000010101100110000110110111100", b"00000000000000000000000000000000"),
	(b"11000010101000000110000111110101", b"01000001000101010101111000111000"), -- 89.5268 + -80.1913 = 9.3355
	(b"11000010100101101110000101110010", b"00000000000000000000000000000000"),
	(b"01000010101001111100101100010100", b"01000001000001110100110100010000"), -- -75.4403 + 83.8966 = 8.45631
	(b"11000001001011100000011100000000", b"00000000000000000000000000000000"),
	(b"11000001100101010000000011111000", b"11000001111011000000010001111000"), -- -10.8767 + -18.6255 = -29.5022
	(b"11000001111110100001011100011000", b"00000000000000000000000000000000"),
	(b"11000010101000110011101001001110", b"11000010111000011100000000010100"), -- -31.2613 + -81.6139 = -112.875
	(b"01000001010010011010101110100000", b"00000000000000000000000000000000"),
	(b"11000001001101001111010000101000", b"00111111101001011011101111000000"), -- 12.6044 + -11.3096 = 1.29479
	(b"01000001001101001001100010111000", b"00000000000000000000000000000000"),
	(b"11000010101011111000010010100110", b"11000010100110001111000110001111"), -- 11.2873 + -87.7591 = -76.4718
	(b"11000001000011001010111111111000", b"00000000000000000000000000000000"),
	(b"11000010011111000001111110000010", b"11000010100011111010010111000000"), -- -8.79296 + -63.0308 = -71.8237
	(b"11000001011000111010110011110000", b"00000000000000000000000000000000"),
	(b"01000010100001110101111001000100", b"01000010010101011101000101001100"), -- -14.2297 + 67.6841 = 53.4544
	(b"11000010010010110010101111111000", b"00000000000000000000000000000000"),
	(b"11000010101000111110000001110000", b"11000011000001001011101100110110"), -- -50.7929 + -81.9384 = -132.731
	(b"11000010101111110000101001001100", b"00000000000000000000000000000000"),
	(b"01000010100100100000001010110110", b"11000001101101000001111001011000"), -- -95.5201 + 73.0053 = -22.5148
	(b"11000010101100100100101000011000", b"00000000000000000000000000000000"),
	(b"11000010000100101101110000011000", b"11000010111110111011100000100100"), -- -89.1447 + -36.7149 = -125.86
	(b"11000010001000010111011101011000", b"00000000000000000000000000000000"),
	(b"11000010000011110000011000100000", b"11000010100110000011111010111100"), -- -40.3665 + -35.756 = -76.1225
	(b"01000010110001100010010110101000", b"00000000000000000000000000000000"),
	(b"01000001010010011110011000011000", b"01000010110111110110001001101011"), -- 99.0735 + 12.6187 = 111.692
	(b"01000001101011110100100111101100", b"00000000000000000000000000000000"),
	(b"11000001000111100001000100110000", b"01000001010000001000001010101000"), -- 21.9111 + -9.8792 = 12.0319
	(b"01000010010101000010001101001011", b"00000000000000000000000000000000"),
	(b"11000010010100111010101110100100", b"00111101111011110100111000000000"), -- 53.0345 + -52.9176 = 0.116848
	(b"01000010010111111011000101011100", b"00000000000000000000000000000000"),
	(b"11000001000100110001010101101000", b"01000010001110101110110000000010"), -- 55.9232 + -9.19273 = 46.7305
	(b"11000010100110001001001101111010", b"00000000000000000000000000000000"),
	(b"11000010100101011011010111001010", b"11000011000101110010010010100010"), -- -76.288 + -74.8551 = -151.143
	(b"01000001010110100001101011111000", b"00000000000000000000000000000000"),
	(b"11000010100101110011001110110010", b"11000010011101111110000010100110"), -- 13.6316 + -75.601 = -61.9694
	(b"11000010101110000100111111100111", b"00000000000000000000000000000000"),
	(b"11000001001101110011100111101000", b"11000010110011110011011100100100"), -- -92.1561 + -11.4516 = -103.608
	(b"01000010011001010111011111101100", b"00000000000000000000000000000000"),
	(b"01000010010110101111111001010100", b"01000010111000000011101100100000"), -- 57.3671 + 54.7484 = 112.115
	(b"11000001110000010111110110111000", b"00000000000000000000000000000000"),
	(b"11000010101000101011000101110010", b"11000010110100110001000011100000"), -- -24.1864 + -81.3466 = -105.533
	(b"01000010011101100011101100101000", b"00000000000000000000000000000000"),
	(b"11000001111100100110110101001100", b"01000001111110100000100100000100"), -- 61.5578 + -30.3034 = 31.2544
	(b"11000010010111110001000000111001", b"00000000000000000000000000000000"),
	(b"11000010000110010101000100100100", b"11000010101111000011000010101110"), -- -55.7658 + -38.3292 = -94.0951
	(b"11000001110100011011010000100000", b"00000000000000000000000000000000"),
	(b"01000001101110001010100010011000", b"11000000010010000101110001000000"), -- -26.213 + 23.0823 = -3.13063
	(b"01000010001101111100110011000000", b"00000000000000000000000000000000"),
	(b"01000000010111010001101101000000", b"01000010010001011001111001110100"), -- 45.95 + 3.45479 = 49.4047
	(b"01000010000100101000000010011111", b"00000000000000000000000000000000"),
	(b"11000001000100110000100110100000", b"01000001110110110111110001101110"), -- 36.6256 + -9.18985 = 27.4358
	(b"11000010101011111110110101110111", b"00000000000000000000000000000000"),
	(b"01000010110001110101000111101000", b"01000001001110110010001110001000"), -- -87.9638 + 99.66 = 11.6962
	(b"11000010010011111010111110010111", b"00000000000000000000000000000000"),
	(b"11000010101011101101100101010110", b"11000011000010110101100010010001"), -- -51.9215 + -87.4245 = -139.346
	(b"11000010100100110001000000001010", b"00000000000000000000000000000000"),
	(b"11000001111001100001100100010000", b"11000010110011001001011001001110"), -- -73.5313 + -28.7622 = -102.294
	(b"01000001100110000110101110000000", b"00000000000000000000000000000000"),
	(b"11000010011010011100011010000100", b"11000010000111011001000011000100"), -- 19.0525 + -58.4439 = -39.3914
	(b"11000010100001101101010101100010", b"00000000000000000000000000000000"),
	(b"11000010010010001111101110100011", b"11000010111010110101001100110100"), -- -67.4168 + -50.2457 = -117.663
	(b"11000001111110111010110110001000", b"00000000000000000000000000000000"),
	(b"11000010001001101100111011001000", b"11000010100100100101001011000110"), -- -31.4597 + -41.7019 = -73.1617
	(b"11000001101011110110010101000100", b"00000000000000000000000000000000"),
	(b"01000001000001010001011100001000", b"11000001010110011011001110000000"), -- -21.9244 + 8.31812 = -13.6063
	(b"01000010100110110011010110011100", b"00000000000000000000000000000000"),
	(b"11000010010101001001101011011000", b"01000001110000111010000011000000"), -- 77.6047 + -53.1512 = 24.4535
	(b"11000010100100010110001011110011", b"00000000000000000000000000000000"),
	(b"11000010100110110000010001000000", b"11000011000101100011001110011010"), -- -72.6933 + -77.5083 = -150.202
	(b"11000010101111100011000110010111", b"00000000000000000000000000000000"),
	(b"11000001111001000111100001111000", b"11000010111101110100111110110101"), -- -95.0969 + -28.5588 = -123.656
	(b"01000001110000100100111010101000", b"00000000000000000000000000000000"),
	(b"11000010101110001010011010111001", b"11000010100010000001001100001111"), -- 24.2884 + -92.3256 = -68.0372
	(b"00111111110110001110000110000000", b"00000000000000000000000000000000"),
	(b"11000010101010110010001101010010", b"11000010101001111011111111001100"), -- 1.69438 + -85.569 = -83.8746
	(b"01000010101010011100000100101010", b"00000000000000000000000000000000"),
	(b"11000010101011100110100110001000", b"11000000000101010000101111000000"), -- 84.8773 + -87.2061 = -2.32884
	(b"01000010000000101010100010011110", b"00000000000000000000000000000000"),
	(b"11000000011111000110101111000000", b"01000001111001011100001111000100"), -- 32.6647 + -3.94408 = 28.7206
	(b"01000010110000110100001101111001", b"00000000000000000000000000000000"),
	(b"01000001100100101110110111010000", b"01000010111001111111111011101101"), -- 97.6318 + 18.3661 = 115.998
	(b"11000010010010001110110100110110", b"00000000000000000000000000000000"),
	(b"11000010100100101011010010101100", b"11000010111101110010101101000111"), -- -50.2317 + -73.3529 = -123.585
	(b"11000010000010001010101100111000", b"00000000000000000000000000000000"),
	(b"11000010100100111000000111001001", b"11000010110101111101011101100101"), -- -34.1672 + -73.7535 = -107.921
	(b"01000000110100010110000000000000", b"00000000000000000000000000000000"),
	(b"11000010101001010001000000011100", b"11000010100101111111101000011100"), -- 6.54297 + -82.5315 = -75.9885
	(b"01000010000100101000000101111010", b"00000000000000000000000000000000"),
	(b"01000010010101110001011111000000", b"01000010101101001100110010011101"), -- 36.6264 + 53.7732 = 90.3996
	(b"01000010100011100110100011100010", b"00000000000000000000000000000000"),
	(b"11000001111110101101001101100000", b"01000010000111110110100000010100"), -- 71.2048 + -31.3532 = 39.8516
	(b"01000001010011000100000000000000", b"00000000000000000000000000000000"),
	(b"01000010001110000101010111101000", b"01000010011010110110010111101000"), -- 12.7656 + 46.0839 = 58.8495
	(b"01000010100101100001101000000010", b"00000000000000000000000000000000"),
	(b"10111111100001111101100101000000", b"01000010100100111111101010011101"), -- 75.0508 + -1.06132 = 73.9895
	(b"01000010001110000010001110110110", b"00000000000000000000000000000000"),
	(b"11000010101100111110001000111100", b"11000010001011111010000011000010"), -- 46.0349 + -89.9419 = -43.907
	(b"11000001010111001111111110011000", b"00000000000000000000000000000000"),
	(b"01000010101001000100010101111110", b"01000010100010001010010110001011"), -- -13.8124 + 82.1357 = 68.3233
	(b"11000010101101001110000111111100", b"00000000000000000000000000000000"),
	(b"10111111011100100100110110000000", b"11000010101101101100011010010111"), -- -90.4414 + -0.946495 = -91.3879
	(b"01000001111101111101011000111100", b"00000000000000000000000000000000"),
	(b"10111111111110000001110110000000", b"01000001111010000101010001100100"), -- 30.9796 + -1.9384 = 29.0412
	(b"11000010101011100110011010111010", b"00000000000000000000000000000000"),
	(b"11000001100101101110011011110100", b"11000010110101000010000001110111"), -- -87.2006 + -18.8628 = -106.063
	(b"01000001101010011010010001100100", b"00000000000000000000000000000000"),
	(b"01000010000111100100010011000100", b"01000010011100110001011011110110"), -- 21.2053 + 39.5672 = 60.7724
	(b"01000010000011011110000101100100", b"00000000000000000000000000000000"),
	(b"01000010000101010011001000010000", b"01000010100100011000100110111010"), -- 35.4701 + 37.2989 = 72.769
	(b"11000010000000100000000101110000", b"00000000000000000000000000000000"),
	(b"11000010001101100010111100111100", b"11000010100111000001100001010110"), -- -32.5014 + -45.5461 = -78.0475
	(b"11000010100111110001111111111100", b"00000000000000000000000000000000"),
	(b"01000010101011001000000011110110", b"01000000110101100000111110100000"), -- -79.5625 + 86.2519 = 6.68941
	(b"01000010101111110000111110100010", b"00000000000000000000000000000000"),
	(b"11000010100101101011011000111010", b"01000001101000010110010110100000"), -- 95.5305 + -75.3559 = 20.1746
	(b"01000010100000111011010100011011", b"00000000000000000000000000000000"),
	(b"11000010100111001111101101011011", b"11000001010010100011001000000000"), -- 65.8537 + -78.4909 = -12.6372
	(b"01000010101100101110011000110100", b"00000000000000000000000000000000"),
	(b"01000010101010110101100011011110", b"01000011001011110001111110001001"), -- 89.4496 + 85.6736 = 175.123
	(b"11000010110001000111111001101011", b"00000000000000000000000000000000"),
	(b"11000010110000011100011110010100", b"11000011010000110010001100000000"), -- -98.2469 + -96.8898 = -195.137
	(b"11000001111011110111011000011000", b"00000000000000000000000000000000"),
	(b"11000010100010100111101110101000", b"11000010110001100101100100101110"), -- -29.9327 + -69.2415 = -99.1742
	(b"11000010110000101111111100111100", b"00000000000000000000000000000000"),
	(b"11000010000010111001100100101000", b"11000011000001000110010111101000"), -- -97.4985 + -34.8996 = -132.398
	(b"01000001100011101001110101001000", b"00000000000000000000000000000000"),
	(b"11000000110110011111111011010000", b"01000001001100000011101100101000"), -- 17.8268 + -6.81236 = 11.0144
	(b"11000001101111111011101000000000", b"00000000000000000000000000000000"),
	(b"01000001111110000111001110001000", b"01000000111000101110011000100000"), -- -23.9658 + 31.0564 = 7.09059
	(b"01000010000010000000111100101100", b"00000000000000000000000000000000"),
	(b"11000010011001100010011010000100", b"11000001101111000010111010110000"), -- 34.0148 + -57.5376 = -23.5228
	(b"11000010001110001011010101001111", b"00000000000000000000000000000000"),
	(b"11000001110001001000101100101000", b"11000010100011010111110101110010"), -- -46.1771 + -24.5679 = -70.745
	(b"01000010010110110110100011111100", b"00000000000000000000000000000000"),
	(b"01000001101110101011111010010000", b"01000010100111000110010000100010"), -- 54.8525 + 23.343 = 78.1956
	(b"11000010101001100001100110100101", b"00000000000000000000000000000000"),
	(b"01000010101011101001110101011110", b"01000000100010000011101110010000"), -- -83.0501 + 87.3074 = 4.25727
	(b"11000001101100001011100100111100", b"00000000000000000000000000000000"),
	(b"10111111111100010010000111000000", b"11000001101111111100101101011000"), -- -22.0904 + -1.88384 = -23.9743
	(b"01000010101000010111100101101100", b"00000000000000000000000000000000"),
	(b"01000010011100101110101011111010", b"01000011000011010111011101110100"), -- 80.7372 + 60.7295 = 141.467
	(b"11000000001111010000111010000000", b"00000000000000000000000000000000"),
	(b"01000000001001010110111001000000", b"10111110101111010000001000000000"), -- -2.95401 + 2.58485 = -0.369156
	(b"01000010100101111001010001010110", b"00000000000000000000000000000000"),
	(b"01000010100000111100010101111000", b"01000011000011011010110011100111"), -- 75.7897 + 65.8857 = 141.675
	(b"01000010000001011111101110100000", b"00000000000000000000000000000000"),
	(b"01000010010011001011000001111000", b"01000010101010010101011000001100"), -- 33.4957 + 51.1723 = 84.6681
	(b"11000001100110011010101111010000", b"00000000000000000000000000000000"),
	(b"11000010101100100000100110011100", b"11000010110110000111010010010000"), -- -19.2089 + -89.0188 = -108.228
	(b"11000010101000100110001001000010", b"00000000000000000000000000000000"),
	(b"01000010101111001100110000011010", b"01000001010100110100111011000000"), -- -81.1919 + 94.3986 = 13.2067
	(b"01000000101101011010110011000000", b"00000000000000000000000000000000"),
	(b"01000000111100001110100010010000", b"01000001010100110100101010101000"), -- 5.67734 + 7.52839 = 13.2057
	(b"11000000000011011000010111000000", b"00000000000000000000000000000000"),
	(b"01000001010010000011010000010000", b"01000001001001001101001010100000"), -- -2.21129 + 12.5127 = 10.3014
	(b"01000010100100001110101010000110", b"00000000000000000000000000000000"),
	(b"01000010000000111000110110111100", b"01000010110100101011000101100100"), -- 72.4581 + 32.8884 = 105.346
	(b"01000001000110011010010010001000", b"00000000000000000000000000000000"),
	(b"01000010110001010011100011000100", b"01000010110110000110110101010101"), -- 9.60267 + 98.6109 = 108.214
	(b"01000010010000010111110100110001", b"00000000000000000000000000000000"),
	(b"10111111010000101001110100000000", b"01000010001111100111001010111101"), -- 48.3723 + -0.760208 = 47.612
	(b"11000010101111110011011000011111", b"00000000000000000000000000000000"),
	(b"01000010001001101010100100110110", b"11000010010101111100001100001000"), -- -95.6057 + 41.6652 = -53.9405
	(b"11000000111010100000111111000000", b"00000000000000000000000000000000"),
	(b"01000001111110101010000111101000", b"01000001110000000001110111111000"), -- -7.31442 + 31.3291 = 24.0146
	(b"01000000110110111001100011010000", b"00000000000000000000000000000000"),
	(b"01000010100011000001100110001110", b"01000010100110011101001100011011"), -- 6.8624 + 70.0499 = 76.9123
	(b"01000010001001111110101000001111", b"00000000000000000000000000000000"),
	(b"01000010100110101011011011110110", b"01000010111011101010101111111110"), -- 41.9786 + 77.3573 = 119.336
	(b"11000001001000001110111011111000", b"00000000000000000000000000000000"),
	(b"11000010100000000111010100001010", b"11000010100101001001001011101001"), -- -10.0583 + -64.2286 = -74.2869
	(b"01000010110000011011100011111111", b"00000000000000000000000000000000"),
	(b"00111111110000010101111100000000", b"01000010110001001011111001111011"), -- 96.8613 + 1.51071 = 98.372
	(b"01000000111111001101011010110000", b"00000000000000000000000000000000"),
	(b"01000001000100100100100110010000", b"01000001100010000101101001110100"), -- 7.90121 + 9.14296 = 17.0442
	(b"11000010100110000010010011110111", b"00000000000000000000000000000000"),
	(b"11000010000101010110101111100000", b"11000010111000101101101011100111"), -- -76.0722 + -37.3553 = -113.428
	(b"01000000000000011010111000100000", b"00000000000000000000000000000000"),
	(b"01000010110000110000100111100110", b"01000010110001110001011101010111"), -- 2.02625 + 97.5193 = 99.5456
	(b"01000001101001011110000011011000", b"00000000000000000000000000000000"),
	(b"11000010100111101001101011000110", b"11000010011010100100010100100000"), -- 20.7348 + -79.3023 = -58.5675
	(b"01000001100000100001010101011000", b"00000000000000000000000000000000"),
	(b"11000001100001011001101111001000", b"10111110111000011001110000000000"), -- 16.2604 + -16.7011 = -0.440643
	(b"11000001100110100100010010110100", b"00000000000000000000000000000000"),
	(b"11000010010110000000001010111111", b"11000010100100101001001010001100"), -- -19.2835 + -54.0027 = -73.2862
	(b"01000010010010100101010110000101", b"00000000000000000000000000000000"),
	(b"11000010011000100010010010011100", b"11000000101111100111100010111000"), -- 50.5835 + -56.5358 = -5.95224
	(b"01000010101110000100101100110001", b"00000000000000000000000000000000"),
	(b"01000001000101110000111110011000", b"01000010110010110010110100100100"), -- 92.1469 + 9.44131 = 101.588
	(b"11000010011001011101000010000000", b"00000000000000000000000000000000"),
	(b"01000010001101111110110011110100", b"11000001001101111000111000110000"), -- -57.4536 + 45.9814 = -11.4722
	(b"01000001110100000011100001001100", b"00000000000000000000000000000000"),
	(b"11000010110001001101011011101100", b"11000010100100001100100011011001"), -- 26.0275 + -98.4198 = -72.3923
	(b"11000010100000011010001010001100", b"00000000000000000000000000000000"),
	(b"11000010010010101000110001111110", b"11000010111001101110100011001011"), -- -64.8175 + -50.6372 = -115.455
	(b"01000010011001011000010101000110", b"00000000000000000000000000000000"),
	(b"01000010000110111001110011100100", b"01000010110000001001000100010101"), -- 57.3801 + 38.9032 = 96.2834
	(b"01000001010101110011011010111000", b"00000000000000000000000000000000"),
	(b"11000001110000001010111111010000", b"11000001001010100010100011101000"), -- 13.4509 + -24.0858 = -10.635
	(b"01000010100110111100000001100110", b"00000000000000000000000000000000"),
	(b"11000010100101001000011010000010", b"01000000011001110011110010000000"), -- 77.8758 + -74.2627 = 3.61307
	(b"01000001101111111110000100100100", b"00000000000000000000000000000000"),
	(b"01000010100111000101100101001110", b"01000010110011000101000110010111"), -- 23.9849 + 78.1744 = 102.159
	(b"01000010100101100100101010001010", b"00000000000000000000000000000000"),
	(b"11000010101010101010000110110010", b"11000001001000101011100101000000"), -- 75.1456 + -85.3158 = -10.1702
	(b"11000010100111010110111101001011", b"00000000000000000000000000000000"),
	(b"11000001110111100001010100010000", b"11000010110101001111010010001111"), -- -78.7174 + -27.7603 = -106.478
	(b"01000010101001000010110011101010", b"00000000000000000000000000000000"),
	(b"01000010010100011011010000110001", b"01000011000001101000001110000001"), -- 82.0877 + 52.426 = 134.514
	(b"01000010010110000010110011000001", b"00000000000000000000000000000000"),
	(b"01000010010011000111010100000000", b"01000010110100100101000011100000"), -- 54.0437 + 51.1143 = 105.158
	(b"11000010000110100011101110101000", b"00000000000000000000000000000000"),
	(b"01000010101110000101111010100011", b"01000010010101101000000110011110"), -- -38.5583 + 92.1848 = 53.6266
	(b"11000001110111001001011000011000", b"00000000000000000000000000000000"),
	(b"11000010101100001010001111011010", b"11000010111001111100100101100000"), -- -27.5733 + -88.32 = -115.893
	(b"01000010010010110111111101111100", b"00000000000000000000000000000000"),
	(b"11000010010101000100100000001001", b"11000000000011001000100011010000"), -- 50.8745 + -53.0703 = -2.19585
	(b"01000010101000010001011100100101", b"00000000000000000000000000000000"),
	(b"11000000101000101110011000110000", b"01000010100101101110100011000010"), -- 80.5452 + -5.0906 = 75.4546
	(b"01000010100011101100101111001101", b"00000000000000000000000000000000"),
	(b"11000000101110100111111001010000", b"01000010100000110010001111101000"), -- 71.398 + -5.82792 = 65.5701
	(b"11000010000001111110011001111000", b"00000000000000000000000000000000"),
	(b"01000010100100010100000110000000", b"01000010000110101001110010001000"), -- -33.9751 + 72.6279 = 38.6529
	(b"01000010100100111010100100011010", b"00000000000000000000000000000000"),
	(b"11000010100010100000000001101001", b"01000000100110101000101100010000"), -- 73.8303 + -69.0008 = 4.82948
	(b"01000010101000010011011001010100", b"00000000000000000000000000000000"),
	(b"11000010100000111101010011010010", b"01000001011010110000110000010000"), -- 80.6061 + -65.9157 = 14.6904
	(b"00111111010010110010101000000000", b"00000000000000000000000000000000"),
	(b"01000010010100100011101010110100", b"01000010010101010110011101011100"), -- 0.79361 + 52.5573 = 53.3509
	(b"01000010011010000110000101011100", b"00000000000000000000000000000000"),
	(b"01000001111100010000111110111000", b"01000010101100000111010010011100"), -- 58.0951 + 30.1327 = 88.2278
	(b"11000010101010010010100111111100", b"00000000000000000000000000000000"),
	(b"01000010100100111110010001100001", b"11000001001010100010110011011000"), -- -84.582 + 73.9461 = -10.6359
	(b"01000010001100000100111000101100", b"00000000000000000000000000000000"),
	(b"11000010100010111000101001000100", b"11000001110011011000110010111000"), -- 44.0763 + -69.7701 = -25.6937
	(b"01000001011100001001011001100000", b"00000000000000000000000000000000"),
	(b"11000010101110000010111001011010", b"11000010100110100001101110001110"), -- 15.0367 + -92.0905 = -77.0538
	(b"11000010000000110110111000111100", b"00000000000000000000000000000000"),
	(b"00111110010000011110000000000000", b"11000010000000101010110001011100"), -- -32.8577 + 0.189331 = -32.6683
	(b"11000010100000100100011010111010", b"00000000000000000000000000000000"),
	(b"11000001110110110111111000110100", b"11000010101110010010011001000111"), -- -65.1381 + -27.4366 = -92.5748
	(b"11000001110110011000111000001100", b"00000000000000000000000000000000"),
	(b"01000000100100111001111011010000", b"11000001101101001010011001011000"), -- -27.1944 + 4.61314 = -22.5812
	(b"01000001011011100110011100000000", b"00000000000000000000000000000000"),
	(b"01000010100111011000010000110100", b"01000010101110110101000100010100"), -- 14.9001 + 78.7582 = 93.6584
	(b"01000010101011100001010100001000", b"00000000000000000000000000000000"),
	(b"01000001111011010001001110010000", b"01000010111010010101100111101100"), -- 87.0411 + 29.6346 = 116.676
	(b"01000010101110101011001010011010", b"00000000000000000000000000000000"),
	(b"11000010011100001010100111100000", b"01000010000001001011101101010100"), -- 93.3488 + -60.1659 = 33.1829
	(b"01000001100001111110100110100100", b"00000000000000000000000000000000"),
	(b"01000010100001111100101000100100", b"01000010101010011100010010001101"), -- 16.9891 + 67.8948 = 84.8839
	(b"11000010010011100110010011010000", b"00000000000000000000000000000000"),
	(b"01000010011000011101110111010111", b"01000000100110111100100000111000"), -- -51.5984 + 56.4666 = 4.86819
	(b"01000010010101111010100001000001", b"00000000000000000000000000000000"),
	(b"11000010011001110101011100000000", b"11000000011110101110101111110000"), -- 53.9143 + -57.835 = -3.92065
	(b"11000010011010100010101100000110", b"00000000000000000000000000000000"),
	(b"01000010000000101101101000101000", b"11000001110011101010000110111100"), -- -58.542 + 32.713 = -25.829
	(b"11000001110100101001101111100100", b"00000000000000000000000000000000"),
	(b"11000010110000111010101111000100", b"11000010111110000101001010111101"), -- -26.3261 + -97.8355 = -124.162
	(b"01000010100010101011101010111110", b"00000000000000000000000000000000"),
	(b"11000010010011000011111101000100", b"01000001100100100110110001110000"), -- 69.3647 + -51.0618 = 18.3029
	(b"01000010110000111011111110011001", b"00000000000000000000000000000000"),
	(b"11000010101101100001100101001111", b"01000000110110100110010010100000"), -- 97.8742 + -91.0494 = 6.82478
	(b"01000010100010000011100110011110", b"00000000000000000000000000000000"),
	(b"11000010011000110000100111000100", b"01000001001101011010010111100000"), -- 68.1125 + -56.7595 = 11.353
	(b"01000001101011010101111110011100", b"00000000000000000000000000000000"),
	(b"11000010100110001110010011101100", b"11000010010110110001101000001010"), -- 21.6717 + -76.4471 = -54.7754
	(b"01000001101001011100001011010100", b"00000000000000000000000000000000"),
	(b"01000010010111110010111000001000", b"01000010100110010000011110111001"), -- 20.7201 + 55.795 = 76.5151
	(b"01000001100100000011010001110000", b"00000000000000000000000000000000"),
	(b"01000010100111101100101010111111", b"01000010110000101101011111011011"), -- 18.0256 + 79.396 = 97.4216
	(b"01000010100010010100010001100001", b"00000000000000000000000000000000"),
	(b"01000010011010000000101101100010", b"01000010111111010100101000010010"), -- 68.6336 + 58.0111 = 126.645
	(b"11000010011011011111111100101000", b"00000000000000000000000000000000"),
	(b"11000010011110001110111010000100", b"11000010111100110111011011010110"), -- -59.4992 + -62.2329 = -121.732
	(b"11000000001111100101001101000000", b"00000000000000000000000000000000"),
	(b"11000010011111110100100100101000", b"11000010100001011001011100101110"), -- -2.97383 + -63.8214 = -66.7953
	(b"01000000010000110101101010000000", b"00000000000000000000000000000000"),
	(b"11000010101110101000101011101101", b"11000010101101000111000000011001"), -- 3.0524 + -93.2713 = -90.2189
	(b"01000001010010011111111110010000", b"00000000000000000000000000000000"),
	(b"01000001100100111001000101100100", b"01000001111110001001000100101100"), -- 12.6249 + 18.446 = 31.0709
	(b"01000010001010010110000110000100", b"00000000000000000000000000000000"),
	(b"11000010010000001011111010111000", b"11000000101110101110100110100000"), -- 42.3452 + -48.1862 = -5.84102
	(b"11000010001111010100001000101101", b"00000000000000000000000000000000"),
	(b"01000010110000001100100001000010", b"01000010010001000100111001010111"), -- -47.3146 + 96.3911 = 49.0765
	(b"01000010101111010111100111101110", b"00000000000000000000000000000000"),
	(b"11000010010011011011100100011000", b"01000010001011010011101011000100"), -- 94.7381 + -51.4308 = 43.3074
	(b"11000001101011100111101101001000", b"00000000000000000000000000000000"),
	(b"01000001011101000111100100101000", b"11000000110100001111101011010000"), -- -21.8102 + 15.2796 = -6.53062
	(b"01000010100110011001110100011000", b"00000000000000000000000000000000"),
	(b"11000010001011010111100100111100", b"01000010000001011100000011110100"), -- 76.8068 + -43.3684 = 33.4384
	(b"01000010100110001010110000011100", b"00000000000000000000000000000000"),
	(b"11000001100011110100000000100000", b"01000010011010011011100000101000"), -- 76.3362 + -17.9063 = 58.4298
	(b"11000010011110101111001000101010", b"00000000000000000000000000000000"),
	(b"11000010010111000110111010111100", b"11000010111010111011000001110011"), -- -62.7365 + -55.1081 = -117.845
	(b"01000010100100010000110000100110", b"00000000000000000000000000000000"),
	(b"01000001110011101001100000000100", b"01000010110001001011001000100111"), -- 72.5237 + 25.8242 = 98.348
	(b"11000010100010101100101010111110", b"00000000000000000000000000000000"),
	(b"01000010011111011000000101111111", b"11000000110000001001111111101000"), -- -69.396 + 63.3765 = -6.01952
	(b"01000010101001001001100101110110", b"00000000000000000000000000000000"),
	(b"01000010101010111001001011000110", b"01000011001010000001011000011110"), -- 82.2997 + 85.7867 = 168.086
	(b"01000010110000100010100101100110", b"00000000000000000000000000000000"),
	(b"11000010011001110101111101101111", b"01000010000111001111001101011101"), -- 97.0809 + -57.8432 = 39.2377
	(b"11000010001101100011011000000100", b"00000000000000000000000000000000"),
	(b"01000010001001010001101110000001", b"11000000100010001101010000011000"), -- -45.5527 + 41.2769 = -4.27589
	(b"01000001111111000010010101000000", b"00000000000000000000000000000000"),
	(b"11000010011100011010010110111100", b"11000001111001110010011000111000"), -- 31.5182 + -60.4118 = -28.8937
	(b"01000010000110100001100111111110", b"00000000000000000000000000000000"),
	(b"01000010001000100010010011010100", b"01000010100111100001111101101001"), -- 38.5254 + 40.536 = 79.0613
	(b"01000010101111101010011011010100", b"00000000000000000000000000000000"),
	(b"11000001111011110010001011000000", b"01000010100000101101111000100100"), -- 95.3258 + -29.892 = 65.4339
	(b"11000010100011110110011100001010", b"00000000000000000000000000000000"),
	(b"11000000101000101101010000000000", b"11000010100110011001010001001010"), -- -71.7012 + -5.08838 = -76.7896
	(b"11000010000101100001111010000000", b"00000000000000000000000000000000"),
	(b"11000010100001000111011110000111", b"11000010110011111000011011000111"), -- -37.5298 + -66.2335 = -103.763
	(b"11000000000000011011111101000000", b"00000000000000000000000000000000"),
	(b"01000010000100110000000000100111", b"01000010000010101110010000110011"), -- -2.0273 + 36.7501 = 34.7229
	(b"01000010010101010100010011001100", b"00000000000000000000000000000000"),
	(b"11000010100011001101011101110010", b"11000001100010001101010000110000"), -- 53.3172 + -70.4208 = -17.1036
	(b"11000010001101110011011110100000", b"00000000000000000000000000000000"),
	(b"11000001001010111000101110010000", b"11000010011000100001101010000100"), -- -45.8043 + -10.7216 = -56.5259
	(b"11000010000011010010000010110100", b"00000000000000000000000000000000"),
	(b"11000010011000001111010111111100", b"11000010101101110000101101011000"), -- -35.2819 + -56.2402 = -91.5222
	(b"11000010010011011110110111000111", b"00000000000000000000000000000000"),
	(b"01000010001101011111010011011100", b"11000000101111111100011101011000"), -- -51.4822 + 45.4891 = -5.99308
	(b"01000010001110100001010000011000", b"00000000000000000000000000000000"),
	(b"11000010010111001110100100000110", b"11000001000010110101001110111000"), -- 46.5196 + -55.2276 = -8.70794
	(b"01000010100011000000001101111100", b"00000000000000000000000000000000"),
	(b"11000010001010010010011001000000", b"01000001110111011100000101110000"), -- 70.0068 + -42.2874 = 27.7195
	(b"11000010011101110010011110100000", b"00000000000000000000000000000000"),
	(b"01000010101010001111111010100000", b"01000001101101011010101101000000"), -- -61.7887 + 84.4973 = 22.7086
	(b"01000000100111000001010110000000", b"00000000000000000000000000000000"),
	(b"11000010100010111100101101100110", b"11000010100000100000101000001110"), -- 4.87762 + -69.8973 = -65.0196
	(b"11000010010001100100111110101100", b"00000000000000000000000000000000"),
	(b"11000010101010100000010101011100", b"11000011000001101001011010011001"), -- -49.5778 + -85.0105 = -134.588
	(b"11000001011100000001111111100000", b"00000000000000000000000000000000"),
	(b"01000001111010011011111101110100", b"01000001011000110101111100001000"), -- -15.0078 + 29.2185 = 14.2107
	(b"01000010101011100000001010100100", b"00000000000000000000000000000000"),
	(b"01000010010101011110100010010111", b"01000011000011000111101101111000"), -- 87.0052 + 53.4771 = 140.482
	(b"11000010101001001110011011110100", b"00000000000000000000000000000000"),
	(b"11000001010111110010100011101000", b"11000010110000001100110000010001"), -- -82.4511 + -13.9475 = -96.3986
	(b"11000001100010011110110100010000", b"00000000000000000000000000000000"),
	(b"01000010011110000001100011000000", b"01000010001100110010001000111000"), -- -17.2408 + 62.0242 = 44.7834
	(b"01000010001001100101011010101100", b"00000000000000000000000000000000"),
	(b"11000001101111110000000000101100", b"01000001100011011010110100101100"), -- 41.5846 + -23.8751 = 17.7096
	(b"01000010010111001110000000010000", b"00000000000000000000000000000000"),
	(b"01000010101010100011111010100001", b"01000011000011000101011101010100"), -- 55.2188 + 85.1223 = 140.341
	(b"11000010100101101001100111110010", b"00000000000000000000000000000000"),
	(b"11000010100110111101101011110010", b"11000011000110010011101001110010"), -- -75.3007 + -77.9276 = -153.228
	(b"01000010000111101101100001000000", b"00000000000000000000000000000000"),
	(b"01000010100101010001110100100100", b"01000010111001001000100101000100"), -- 39.7112 + 74.5569 = 114.268
	(b"11000010000101010111010111000100", b"00000000000000000000000000000000"),
	(b"01000010101111011010011001010000", b"01000010011001011101011011011100"), -- -37.365 + 94.8248 = 57.4598
	(b"11000010100101111110001011101000", b"00000000000000000000000000000000"),
	(b"01000001010111011111001011010000", b"11000010011110000100100100011100"), -- -75.9432 + 13.8718 = -62.0714
	(b"11000010001001110101011000101111", b"00000000000000000000000000000000"),
	(b"11000010001111100001010010011111", b"11000010101100101011010101100111"), -- -41.8342 + -47.5201 = -89.3543
	(b"01000010100011110011101000000110", b"00000000000000000000000000000000"),
	(b"01000010001110101110100111000000", b"01000010111011001010111011100110"), -- 71.6133 + 46.7283 = 118.342
	(b"11000010011001110110101011111010", b"00000000000000000000000000000000"),
	(b"11000010100011100110010101001110", b"11000011000000010000110101100110"), -- -57.8545 + -71.1979 = -129.052
	(b"01000010011110111100100111011000", b"00000000000000000000000000000000"),
	(b"01000001111101100100011011110100", b"01000010101110110111011010101001"), -- 62.9471 + 30.7846 = 93.7318
	(b"11000010101110111111011110110110", b"00000000000000000000000000000000"),
	(b"01000010100100001011011100011100", b"11000001101011010000001001101000"), -- -93.9838 + 72.3576 = -21.6262
	(b"11000010101010100010110110010000", b"00000000000000000000000000000000"),
	(b"01000010011111001000011111101100", b"11000001101011111010011001101000"), -- -85.089 + 63.1327 = -21.9563
	(b"01000001111100100000001011010000", b"00000000000000000000000000000000"),
	(b"11000010001010011000010011011100", b"11000001010000100000110111010000"), -- 30.2514 + -42.3797 = -12.1284
	(b"01000010010110001010011011111000", b"00000000000000000000000000000000"),
	(b"01000010100011111111110011110110", b"01000010111111000101000001110010"), -- 54.1631 + 71.9941 = 126.157
	(b"01000010001111000010111101000101", b"00000000000000000000000000000000"),
	(b"01000000110001011010001100110000", b"01000010010101001110001110101011"), -- 47.0462 + 6.17617 = 53.2223
	(b"11000010000110001000111110100100", b"00000000000000000000000000000000"),
	(b"11000010011100111110011000101000", b"11000010110001100011101011100110"), -- -38.1403 + -60.9748 = -99.115
	(b"01000010011000000011011010001100", b"00000000000000000000000000000000"),
	(b"11000010101100110001001110100011", b"11000010000001011111000010111010"), -- 56.0533 + -89.5384 = -33.4851
	(b"11000001101101110000100111011000", b"00000000000000000000000000000000"),
	(b"11000001111101000111011011000000", b"11000010010101011100000001001100"), -- -22.8798 + -30.558 = -53.4378
	(b"01000001100011111011110001010100", b"00000000000000000000000000000000"),
	(b"01000010100110110010001111100111", b"01000010101111110001001011111100"), -- 17.967 + 77.5701 = 95.5371
	(b"01000000110110000110011110110000", b"00000000000000000000000000000000"),
	(b"11000010011110011001000110100100", b"11000010010111101000010010101110"), -- 6.76266 + -62.3922 = -55.6296
	(b"11000010100010011101010001011000", b"00000000000000000000000000000000"),
	(b"11000000000001011110010111000000", b"11000010100011100000001110000110"), -- -68.9147 + -2.09215 = -71.0069
	(b"01000010100101011100011110011000", b"00000000000000000000000000000000"),
	(b"11000010000100111100011100111000", b"01000010000101111100011111111000"), -- 74.8898 + -36.9445 = 37.9453
	(b"11000010101010101000110100000100", b"00000000000000000000000000000000"),
	(b"01000010010001010000100001001100", b"11000010000100000001000110111100"), -- -85.2754 + 49.2581 = -36.0173
	(b"11000010011001001001010110010000", b"00000000000000000000000000000000"),
	(b"11000010110000001000111110110011", b"11000011000110010110110100111110"), -- -57.1461 + -96.2807 = -153.427
	(b"01000001011011111000101010011000", b"00000000000000000000000000000000"),
	(b"01000010011011000011000111110000", b"01000010100101000000101001001011"), -- 14.9713 + 59.0488 = 74.0201
	(b"01000010001001001011010101101000", b"00000000000000000000000000000000"),
	(b"01000010100111010010110111011100", b"01000010111011111000100010010000"), -- 41.1772 + 78.5896 = 119.767
	(b"11000001101010101100010110011100", b"00000000000000000000000000000000"),
	(b"11000010100001011011010101011000", b"11000010101100000110011010111111"), -- -21.3465 + -66.8542 = -88.2007
	(b"01000010110001100101011000111000", b"00000000000000000000000000000000"),
	(b"11000001100011101101110010101000", b"01000010101000101001111100001110"), -- 99.1684 + -17.8577 = 81.3107
	(b"11000010100001110100011010101001", b"00000000000000000000000000000000"),
	(b"01000010001111101001011001110011", b"11000001100111111110110110111110"), -- -67.638 + 47.6469 = -19.9911
	(b"11000010101000101001011100011000", b"00000000000000000000000000000000"),
	(b"11000010100100011101011010011010", b"11000011000110100011011011011001"), -- -81.2951 + -72.9191 = -154.214
	(b"01000010101011100001110010101001", b"00000000000000000000000000000000"),
	(b"11000010100011000001100101110101", b"01000001100010000000110011010000"), -- 87.056 + -70.0497 = 17.0063
	(b"01000010100111000111110100011110", b"00000000000000000000000000000000"),
	(b"01000001111110111001101100011000", b"01000010110110110110001111100100"), -- 78.2444 + 31.4507 = 109.695
	(b"01000010001011011010110111000000", b"00000000000000000000000000000000"),
	(b"01000010000111100100011110110001", b"01000010101001011111101010111000"), -- 43.4197 + 39.57 = 82.9897
	(b"11000010100001100100111001001000", b"00000000000000000000000000000000"),
	(b"11000001100011110001111010000000", b"11000010101010100001010111101000"), -- -67.1529 + -17.8899 = -85.0428
	(b"11000010000000100101101110011100", b"00000000000000000000000000000000"),
	(b"11000000100101110110011011100000", b"11000010000101010100100001111000"), -- -32.5895 + -4.73131 = -37.3208
	(b"01000010001011111001011000011001", b"00000000000000000000000000000000"),
	(b"11000001100101010011000000000100", b"01000001110010011111110000101110"), -- 43.8966 + -18.6484 = 25.2481
	(b"01000001010101100001010110001000", b"00000000000000000000000000000000"),
	(b"01000010100000000011111111011110", b"01000010100110110000001010001111"), -- 13.3803 + 64.1247 = 77.505
	(b"11000001100011011000111111000100", b"00000000000000000000000000000000"),
	(b"11000010001000101000001001011100", b"11000010011010010100101000111110"), -- -17.6952 + -40.6273 = -58.3225
	(b"01000010101101110010111011001011", b"00000000000000000000000000000000"),
	(b"01000010010100101101111111010100", b"01000011000100000100111101011010"), -- 91.5914 + 52.7186 = 144.31
	(b"11000010101000010101101100001100", b"00000000000000000000000000000000"),
	(b"01000010100101001010110001011011", b"11000000110010101110101100010000"), -- -80.6778 + 74.3366 = -6.34119
	(b"11000010000010111011010000111000", b"00000000000000000000000000000000"),
	(b"11000010001011101101100001001010", b"11000010100111010100011001000001"), -- -34.926 + -43.7112 = -78.6372
	(b"01000010101001011001001011111010", b"00000000000000000000000000000000"),
	(b"11000010100000010110011101101110", b"01000001100100001010111000110000"), -- 82.7871 + -64.702 = 18.0851
	(b"01000010000100010001100001011111", b"00000000000000000000000000000000"),
	(b"01000010001011010110000110110000", b"01000010100111110011110100001000"), -- 36.2738 + 43.3454 = 79.6192
	(b"11000010010111011010111111101100", b"00000000000000000000000000000000"),
	(b"01000010001100110100011100100000", b"11000001001010011010001100110000"), -- -55.4218 + 44.8195 = -10.6023
	(b"01000010101000001011001100101010", b"00000000000000000000000000000000"),
	(b"01000001100100110010111001001100", b"01000010110001010111111010111101"), -- 80.3499 + 18.3976 = 98.7475
	(b"11000010101100100000011010010110", b"00000000000000000000000000000000"),
	(b"01000000101001110011011110110000", b"11000010101001111001001100011011"), -- -89.0129 + 5.22555 = -83.7873
	(b"01000001100100001110000000010000", b"00000000000000000000000000000000"),
	(b"11000010110001001111100000010001", b"11000010101000001100000000001101"), -- 18.1094 + -98.4845 = -80.3751
	(b"01000010101011000011011001100011", b"00000000000000000000000000000000"),
	(b"01000010100111100010011000010011", b"01000011001001010010111000111011"), -- 86.1062 + 79.0744 = 165.181
	(b"11000010110000000010100000010000", b"00000000000000000000000000000000"),
	(b"01000010110000110011100101001000", b"00111111110001000100111000000000"), -- -96.0782 + 97.6119 = 1.53363
	(b"11000001110100100101000110110100", b"00000000000000000000000000000000"),
	(b"01000010011101010000000101110111", b"01000010000010111101100010011101"), -- -26.2899 + 61.2514 = 34.9615
	(b"01000000110111100001110111010000", b"00000000000000000000000000000000"),
	(b"11000001110011001110111110000000", b"11000001100101010110100000001100"), -- 6.94114 + -25.6169 = -18.6758
	(b"01000010001111110110100010010110", b"00000000000000000000000000000000"),
	(b"10111110100011110101000100000000", b"01000010001111100100100111110100"), -- 47.8521 + -0.279915 = 47.5722
	(b"01000010011111110000110100101100", b"00000000000000000000000000000000"),
	(b"11000010101111111001101001011110", b"11000010000000000010011110010000"), -- 63.7629 + -95.8015 = -32.0386
	(b"01000010010110100011000011001000", b"00000000000000000000000000000000"),
	(b"11000010001100110111011000011111", b"01000001000110101110101010100100"), -- 54.5476 + -44.8654 = 9.68229
	(b"01000001000011010001010011110000", b"00000000000000000000000000000000"),
	(b"01000010100011011110111011000110", b"01000010100111111001000101100100"), -- 8.81761 + 70.9664 = 79.784
	(b"01000010100010111110111001011000", b"00000000000000000000000000000000"),
	(b"11000010100100100001011001000010", b"11000000010001001111110101000000"), -- 69.9655 + -73.0435 = -3.07796
	(b"01000010101100001101110110100110", b"00000000000000000000000000000000"),
	(b"01000010100100000011111111000111", b"01000011001000001000111010110110"), -- 88.4329 + 72.1246 = 160.557
	(b"11000001110010110111000000111100", b"00000000000000000000000000000000"),
	(b"11000010101010111111010110010110", b"11000010110111101101000110100101"), -- -25.4298 + -85.9797 = -111.409
	(b"01000001010001110011001011001000", b"00000000000000000000000000000000"),
	(b"11000001111111111110011011001000", b"11000001100111000100110101100100"), -- 12.4499 + -31.9877 = -19.5378
	(b"11000010010101110001100111101100", b"00000000000000000000000000000000"),
	(b"11000010010010000011101111110100", b"11000010110011111010101011110000"), -- -53.7753 + -50.0585 = -103.834
	(b"11000010100110001111000000011000", b"00000000000000000000000000000000"),
	(b"01000010010011111010000101111100", b"11000001110001000111110101101000"), -- -76.4689 + 51.9077 = -24.5612
	(b"01000010101110010100011101101000", b"00000000000000000000000000000000"),
	(b"11000010000110000010101011101110", b"01000010010110100110001111100010"), -- 92.6395 + -38.0419 = 54.5975
	(b"01000010000101110101001101110010", b"00000000000000000000000000000000"),
	(b"11000010011111001110011011100100", b"11000001110010110010011011100100"), -- 37.8315 + -63.2255 = -25.394
	(b"01000010100011111011011010101110", b"00000000000000000000000000000000"),
	(b"11000010001000100110110000111100", b"01000001111110100000001001000000"), -- 71.8568 + -40.6057 = 31.2511
	(b"11000010000101111000001100010100", b"00000000000000000000000000000000"),
	(b"01000010001011100111111100011000", b"01000000101101111110000000100000"), -- -37.878 + 43.6241 = 5.74611
	(b"01000001110000010111001110110100", b"00000000000000000000000000000000"),
	(b"11000001110010100011000000010100", b"10111111100010111100011000000000"), -- 24.1815 + -25.2735 = -1.09198
	(b"11000010100001101111110001101100", b"00000000000000000000000000000000"),
	(b"11000010000010010100101101011000", b"11000010110010111010001000011000"), -- -67.493 + -34.3236 = -101.817
	(b"11000001101001110100100111000000", b"00000000000000000000000000000000"),
	(b"01000010100001011100010101110111", b"01000010001101111110011000001110"), -- -20.911 + 66.8857 = 45.9747
	(b"11000010011101000000100010010100", b"00000000000000000000000000000000"),
	(b"11000010100101101111100010000010", b"11000011000010000111111001100110"), -- -61.0084 + -75.4854 = -136.494
	(b"01000010101010011011010000011010", b"00000000000000000000000000000000"),
	(b"11000010100010000010111110110010", b"01000001100001100001000110100000"), -- 84.8518 + -68.0932 = 16.7586
	(b"01000010001010110100111001110011", b"00000000000000000000000000000000"),
	(b"01000010100101010111110111111100", b"01000010111010110010010100110110"), -- 42.8266 + 74.7461 = 117.573
	(b"11000010101010000111011010000010", b"00000000000000000000000000000000"),
	(b"11000010000100010100010000010000", b"11000010111100010001100010001010"), -- -84.2315 + -36.3165 = -120.548
	(b"01000010001010001011101111101011", b"00000000000000000000000000000000"),
	(b"01000001110101001001101001001100", b"01000010100010011000010010001000"), -- 42.1835 + 26.5753 = 68.7589
	(b"01000001101100101110000011100100", b"00000000000000000000000000000000"),
	(b"01000010101000111111000011111000", b"01000010110100001010100100110001"), -- 22.3598 + 81.9706 = 104.33
	(b"01000010101010101101100100000100", b"00000000000000000000000000000000"),
	(b"01000010101111011011100101010110", b"01000011001101000100100100101101"), -- 85.4239 + 94.862 = 180.286
	(b"11000010101100011001111010111110", b"00000000000000000000000000000000"),
	(b"11000010101111001001101111110111", b"11000011001101110001110101011010"), -- -88.81 + -94.3046 = -183.115
	(b"11000010100101010100001111111100", b"00000000000000000000000000000000"),
	(b"11000010001000010100000010111101", b"11000010111001011110010001011010"), -- -74.6328 + -40.3132 = -114.946
	(b"11000010000011110100110111001100", b"00000000000000000000000000000000"),
	(b"01000010101011011110000000010011", b"01000010010011000111001001011010"), -- -35.826 + 86.9376 = 51.1117
	(b"01000010101110011001100011000010", b"00000000000000000000000000000000"),
	(b"11000010101100100000110100110110", b"01000000011100010111000110000000"), -- 92.7984 + -89.0258 = 3.77255
	(b"01000010010100001111111110011000", b"00000000000000000000000000000000"),
	(b"11000001011011001000011011011000", b"01000010000101011101110111100010"), -- 52.2496 + -14.7829 = 37.4667
	(b"01000010100001000011101011110100", b"00000000000000000000000000000000"),
	(b"00111111101010100111111100000000", b"01000010100001101110010011110000"), -- 66.1151 + 1.332 = 67.4471
	(b"11000010100100011100001111110011", b"00000000000000000000000000000000"),
	(b"11000010011000010001100011011100", b"11000011000000010010100000110000"), -- -72.8827 + -56.2743 = -129.157
	(b"01000010011000000001110000000000", b"00000000000000000000000000000000"),
	(b"01000000110011101110110011100000", b"01000010011110011111100110011100"), -- 56.0273 + 6.46642 = 62.4938
	(b"01000010101100101011100010001010", b"00000000000000000000000000000000"),
	(b"01000001111010101100010101010000", b"01000010111011010110100111011110"), -- 89.3604 + 29.3463 = 118.707
	(b"11000001111101000001001001110000", b"00000000000000000000000000000000"),
	(b"11000010101010111101101100111110", b"11000010111010001101111111011010"), -- -30.509 + -85.9282 = -116.437
	(b"11000010000100011010111111001000", b"00000000000000000000000000000000"),
	(b"01000010100101111110011000000110", b"01000010000111100001110001000100"), -- -36.4217 + 75.9493 = 39.5276
	(b"11000000001010010000100010100000", b"00000000000000000000000000000000"),
	(b"01000010011111111000001011100010", b"01000010011101001111001001011000"), -- -2.64115 + 63.8778 = 61.2367
	(b"11000010100000111111100100010110", b"00000000000000000000000000000000"),
	(b"01000001110111110110100101110000", b"11000010000110000011110101110100"), -- -65.9865 + 27.9265 = -38.06
	(b"11000010100011000111110011011010", b"00000000000000000000000000000000"),
	(b"01000010110001110101000111011110", b"01000001111010110101010000010000"), -- -70.2439 + 99.6599 = 29.416
	(b"11000010100011000001010011011001", b"00000000000000000000000000000000"),
	(b"01000010000101111011011001111100", b"11000010000000000111001100110110"), -- -70.0407 + 37.9282 = -32.1125
	(b"10111111011000110011000110000000", b"00000000000000000000000000000000"),
	(b"11000000001000110110101010100000", b"11000000010111000011011100000000"), -- -0.887474 + -2.55338 = -3.44086
	(b"10111111100111001111001000000000", b"00000000000000000000000000000000"),
	(b"10111111100000101100001110000000", b"11000000000011111101101011000000"), -- -1.22614 + -1.02159 = -2.24773
	(b"11000001111011000011010100001000", b"00000000000000000000000000000000"),
	(b"01000010101010001011001101101110", b"01000010010110110100110001011000"), -- -29.5259 + 84.3504 = 54.8246
	(b"01000000100110111010011011100000", b"00000000000000000000000000000000"),
	(b"01000010100010001011111011001100", b"01000010100100100111100100111010"), -- 4.86412 + 68.3727 = 73.2368
	(b"01000010101101000001011101111010", b"00000000000000000000000000000000"),
	(b"01000010011111110110011100110101", b"01000011000110011110010110001010"), -- 90.0459 + 63.8508 = 153.897
	(b"11000010100011011000110101010011", b"00000000000000000000000000000000"),
	(b"01000001111000111111110101111000", b"11000010001010010001101111101010"), -- -70.776 + 28.4988 = -42.2773
	(b"01000010011001110010010100011010", b"00000000000000000000000000000000"),
	(b"01000000111110100111000101010000", b"01000010100000110011100110100010"), -- 57.7862 + 7.82633 = 65.6126
	(b"01000010001111011001010101110110", b"00000000000000000000000000000000"),
	(b"01000010011100011000011000010000", b"01000010110101111000110111000011"), -- 47.396 + 60.3809 = 107.777
	(b"11000001100010010000000001010000", b"00000000000000000000000000000000"),
	(b"11000010100010010000001100000101", b"11000010101010110100001100011001"), -- -17.1252 + -68.5059 = -85.6311
	(b"11000010011001100111110001100000", b"00000000000000000000000000000000"),
	(b"01000010011010010101011000011100", b"00111111001101100110111100000000"), -- -57.6215 + 58.3341 = 0.712631
	(b"01000010100010001110011111111110", b"00000000000000000000000000000000"),
	(b"01000010101000110000100111000011", b"01000011000101011111100011100000"), -- 68.4531 + 81.5191 = 149.972
	(b"11000010001010011011010110001000", b"00000000000000000000000000000000"),
	(b"01000010011110011001011111000000", b"01000001100111111100010001110000"), -- -42.4273 + 62.3982 = 19.9709
	(b"11000010011100010001001110110100", b"00000000000000000000000000000000"),
	(b"01000010101111101010100101100111", b"01000010000011000011111100011010"), -- -60.2692 + 95.3309 = 35.0616
	(b"11000010000110100110110000100100", b"00000000000000000000000000000000"),
	(b"11000000110010001101011111010000", b"11000010001100111000011100011110"), -- -38.6056 + -6.27634 = -44.882
	(b"01000001100010011010101010001000", b"00000000000000000000000000000000"),
	(b"01000010100001110110101011011010", b"01000010101010011101010101111100"), -- 17.2083 + 67.7087 = 84.917
	(b"01000010010100100110001010011011", b"00000000000000000000000000000000"),
	(b"01000010000010001011111101011010", b"01000010101011011001000011111010"), -- 52.5963 + 34.1869 = 86.7832
	(b"01000010101011000101011010101111", b"00000000000000000000000000000000"),
	(b"01000010100000000101101010100000", b"01000011000101100101100010101000"), -- 86.1693 + 64.177 = 150.346
	(b"01000010001001101100010100011100", b"00000000000000000000000000000000"),
	(b"11000001111001100100110100101000", b"01000001010011100111101000100000"), -- 41.6925 + -28.7877 = 12.9048
	(b"11000010100100000000000010010011", b"00000000000000000000000000000000"),
	(b"01000001100001101100110111011100", b"11000010010111001001101000111000"), -- -72.0011 + 16.8505 = -55.1506
	(b"01000010011000010011001011110100", b"00000000000000000000000000000000"),
	(b"01000001010011011110000100100000", b"01000010100010100101010110011110"), -- 56.2998 + 12.8675 = 69.1672
	(b"01000010001000111001011100001100", b"00000000000000000000000000000000"),
	(b"11000010000101101110100011000000", b"01000000010010101110010011000000"), -- 40.8975 + -37.7273 = 3.17021
	(b"11000001101100110001101000110000", b"00000000000000000000000000000000"),
	(b"11000001110000000000110000010000", b"11000010001110011001001100100000"), -- -22.3878 + -24.0059 = -46.3937
	(b"11000001011010110111110100000000", b"00000000000000000000000000000000"),
	(b"01000010100001100011001010001010", b"01000010010100011000010111010100"), -- -14.718 + 67.0987 = 52.3807
	(b"11000010100010000100011001110010", b"00000000000000000000000000000000"),
	(b"11000001110011101110101001001000", b"11000010101111000000000100000100"), -- -68.1376 + -25.8644 = -94.002
	(b"11000001110000001011000001111100", b"00000000000000000000000000000000"),
	(b"11000010101101101111000000001101", b"11000010111001110001110000101100"), -- -24.0862 + -91.4688 = -115.555
	(b"01000010010110011000010100001000", b"00000000000000000000000000000000"),
	(b"11000010100111010110100111100110", b"11000001110000101001110110001000"), -- 54.3799 + -78.7068 = -24.3269
	(b"01000010101000010011111110010010", b"00000000000000000000000000000000"),
	(b"01000010101000000100100001011010", b"01000011001000001100001111110110"), -- 80.6242 + 80.1413 = 160.765
	(b"01000001000011100011100110001000", b"00000000000000000000000000000000"),
	(b"01000010001110000000010110100100", b"01000010010110111001010000000110"), -- 8.88905 + 46.0055 = 54.8946
	(b"01000001100100010100101101101000", b"00000000000000000000000000000000"),
	(b"11000001111010100111010100010100", b"11000001001100100101001101011000"), -- 18.1618 + -29.3072 = -11.1453
	(b"01000010100011100001100010001010", b"00000000000000000000000000000000"),
	(b"11000010110000000011110000100000", b"11000001110010001000111001011000"), -- 71.0479 + -96.1174 = -25.0695
	(b"01000010010100010101101101011100", b"00000000000000000000000000000000"),
	(b"01000010000111111100001011010100", b"01000010101110001000111100011000"), -- 52.3392 + 39.9403 = 92.2795
	(b"11000010000111001100101100110100", b"00000000000000000000000000000000"),
	(b"01000010000010100111110000101110", b"11000000100100100111100000110000"), -- -39.1984 + 34.6213 = -4.57717
	(b"01000010010100101011010011110010", b"00000000000000000000000000000000"),
	(b"01000010101001110101100010110100", b"01000011000010000101100110010110"), -- 52.6767 + 83.6732 = 136.35
	(b"01000010100011001100100000001110", b"00000000000000000000000000000000"),
	(b"01000001000111011111110100110000", b"01000010101000001000011110110100"), -- 70.3907 + 9.87431 = 80.265
	(b"01000000110101110000101111000000", b"00000000000000000000000000000000"),
	(b"01000010100111100000011101110100", b"01000010101010110111100000110000"), -- 6.72018 + 79.0146 = 85.7347
	(b"11000010001000110111110100001001", b"00000000000000000000000000000000"),
	(b"11000010101111110000011111101110", b"11000011000010000110001100111001"), -- -40.8721 + -95.5155 = -136.388
	(b"11000001000111111101011110110000", b"00000000000000000000000000000000"),
	(b"11000010000001000110111001110010", b"11000010001011000110010001011110"), -- -9.99016 + -33.1079 = -43.098
	(b"11000001011011101110001000111000", b"00000000000000000000000000000000"),
	(b"11000000101100101010010011110000", b"11000001101001000001101001011000"), -- -14.9302 + -5.58263 = -20.5129
	(b"01000001100000001011100110101000", b"00000000000000000000000000000000"),
	(b"11000001111101101100010000100000", b"11000001011011000001010011110000"), -- 16.0907 + -30.8458 = -14.7551
	(b"11000001010100000011101001101000", b"00000000000000000000000000000000"),
	(b"11000001110010110001111110010000", b"11000010000110011001111001100010"), -- -13.0143 + -25.3904 = -38.4047
	(b"01000010011001111000011100000100", b"00000000000000000000000000000000"),
	(b"01000001111000111000100101011000", b"01000010101011001010010111011000"), -- 57.8819 + 28.4421 = 86.3239
	(b"01000010011011001101011111010000", b"00000000000000000000000000000000"),
	(b"01000010100000101111000010000010", b"01000010111110010101110001101010"), -- 59.2108 + 65.4697 = 124.68
	(b"11000010101100000111101111011110", b"00000000000000000000000000000000"),
	(b"01000001111001001011111101111100", b"11000010011011101001011111111110"), -- -88.2419 + 28.5935 = -59.6484
	(b"11000010101111111010100100000100", b"00000000000000000000000000000000"),
	(b"01000001000011000101111001101000", b"11000010101011100001110100110111"), -- -95.8301 + 8.77305 = -87.0571
	(b"01000000111011000110000001010000", b"00000000000000000000000000000000"),
	(b"11000001101101011101111101111000", b"11000001011101011000111011001000"), -- 7.38676 + -22.7341 = -15.3474
	(b"11000001100010010110110011101000", b"00000000000000000000000000000000"),
	(b"11000001100011110001001101010000", b"11000010000011000100000000011100"), -- -17.1782 + -17.8844 = -35.0626
	(b"01000010011100111101010101001111", b"00000000000000000000000000000000"),
	(b"11000000101001011011110001000000", b"01000010010111110001110111000111"), -- 60.9583 + -5.17923 = 55.7791
	(b"01000010100101100100100001000000", b"00000000000000000000000000000000"),
	(b"11000010100011001110011011100000", b"01000000100101100001011000000000"), -- 75.1411 + -70.4509 = 4.69019
	(b"01000001101010100000111101111000", b"00000000000000000000000000000000"),
	(b"00111111101110010001100110000000", b"01000001101101011010000100010000"), -- 21.2576 + 1.44609 = 22.7036
	(b"01000010100000000101110111110100", b"00000000000000000000000000000000"),
	(b"01000010101111110100000000110000", b"01000011000111111100111100010010"), -- 64.1835 + 95.6254 = 159.809
	(b"01000001010000011001000111000000", b"00000000000000000000000000000000"),
	(b"11000010001101000101001010001000", b"11000010000000111110111000011000"), -- 12.0981 + -45.0806 = -32.9825
	(b"11000010011010000011110001110111", b"00000000000000000000000000000000"),
	(b"01000010000111001001010110010100", b"11000001100101110100110111000110"), -- -58.059 + 39.1461 = -18.913
	(b"11000010000011010001010101010100", b"00000000000000000000000000000000"),
	(b"01000010010000001001101001100100", b"01000001010011100001010001000000"), -- -35.2708 + 48.1508 = 12.8799
	(b"11000010001001000111100110011010", b"00000000000000000000000000000000"),
	(b"11000010110001011100010111001000", b"11000011000011000000000101001010"), -- -41.1188 + -98.8863 = -140.005
	(b"01000010101001101011001010110100", b"00000000000000000000000000000000"),
	(b"01000001111100011000100101000000", b"01000010111000110001010100000100"), -- 83.349 + 30.192 = 113.541
	(b"11000001110001000000101100101100", b"00000000000000000000000000000000"),
	(b"11000010011001111001001010001100", b"11000010101001001100110000010001"), -- -24.5055 + -57.8931 = -82.3986
	(b"01000001101011000100111101001100", b"00000000000000000000000000000000"),
	(b"01000001001100111101011111001000", b"01000010000000110001110110011000"), -- 21.5387 + 11.2402 = 32.7789
	(b"01000000100101100101000100010000", b"00000000000000000000000000000000"),
	(b"01000010101001110101110001000010", b"01000010101100001100000101010011"), -- 4.6974 + 83.6802 = 88.3776
	(b"01000001011001011111011100100000", b"00000000000000000000000000000000"),
	(b"01000010010001111101000110110011", b"01000010100000001010011110111110"), -- 14.3728 + 49.9548 = 64.3276
	(b"11000010001011001101111100001100", b"00000000000000000000000000000000"),
	(b"11000010010111101000010111100000", b"11000010110001011011001001110110"), -- -43.2178 + -55.6307 = -98.8486
	(b"01000010100111101011000111100100", b"00000000000000000000000000000000"),
	(b"11000010110000010001000010001000", b"11000001100010010111101010010000"), -- 79.3474 + -96.5323 = -17.1848
	(b"11000000110101110010001010100000", b"00000000000000000000000000000000"),
	(b"11000001110001111011111101101000", b"11000001111111011000100000010000"), -- -6.72298 + -24.9685 = -31.6914
	(b"01000010101001010100001011110110", b"00000000000000000000000000000000"),
	(b"01000010100010000011010111000100", b"01000011000101101011110001011101"), -- 82.6308 + 68.105 = 150.736
	(b"00111111001000100101001110000000", b"00000000000000000000000000000000"),
	(b"01000010010110101111010111011100", b"01000010010111010111111100101010"), -- 0.634087 + 54.7401 = 55.3742
	(b"01000010101111110100111010111010", b"00000000000000000000000000000000"),
	(b"11000010100100011000000000101011", b"01000001101101110011101000111100"), -- 95.6538 + -72.7503 = 22.9034
	(b"01000010010010111011000011100100", b"00000000000000000000000000000000"),
	(b"11000010010000010011001101000010", b"01000000001001111101101000100000"), -- 50.9227 + -48.3001 = 2.62269
	(b"01000000100101001001000101000000", b"00000000000000000000000000000000"),
	(b"11000001111000000000100011111000", b"11000001101110101110010010101000"), -- 4.64273 + -28.0044 = -23.3616
	(b"00111111111110011111010000000000", b"00000000000000000000000000000000"),
	(b"11000010100110000110101100101110", b"11000010100101001000001101011110"), -- 1.95276 + -76.2093 = -74.2566
	(b"01000010100101100010111011110110", b"00000000000000000000000000000000"),
	(b"01000001111101100010110100000000", b"01000010110100111011101000110110"), -- 75.0917 + 30.772 = 105.864
	(b"01000010000010111011011111010100", b"00000000000000000000000000000000"),
	(b"01000001011111101001100010111000", b"01000010010010110101111000000010"), -- 34.9295 + 15.9123 = 50.8418
	(b"01000010011000110111001001111011", b"00000000000000000000000000000000"),
	(b"11000010000101000110000110001100", b"01000001100111100010000111011110"), -- 56.8618 + -37.0953 = 19.7665
	(b"11000010001101111010101110001100", b"00000000000000000000000000000000"),
	(b"11000010100110111000111001110000", b"11000010111101110110010000110110"), -- -45.9175 + -77.7782 = -123.696
	(b"11000010100010000101111101001010", b"00000000000000000000000000000000"),
	(b"11000010011111010100010110110000", b"11000011000000111000000100010001"), -- -68.1861 + -63.3181 = -131.504
	(b"11000010110000000011010010110111", b"00000000000000000000000000000000"),
	(b"11000001100001101001010010101000", b"11000010111000011101100111100001"), -- -96.103 + -16.8226 = -112.926
	(b"11000010100101010100011111010110", b"00000000000000000000000000000000"),
	(b"11000010110001010010110010101000", b"11000011001011010011101000111111"), -- -74.6403 + -98.5872 = -173.228
	(b"11000001100100001001000010010000", b"00000000000000000000000000000000"),
	(b"01000010110001001011000101100000", b"01000010101000001000110100111100"), -- -18.0706 + 98.3464 = 80.2758
	(b"11000010101000011110110100011100", b"00000000000000000000000000000000"),
	(b"01000010010000100110010100001100", b"11000010000000010111010100101100"), -- -80.9631 + 48.5987 = -32.3644
	(b"01000010100010111101010110100100", b"00000000000000000000000000000000"),
	(b"11000010101000000001101011101010", b"11000001001000100010101000110000"), -- 69.9173 + -80.0526 = -10.1353
	(b"01000010001110111110011111001100", b"00000000000000000000000000000000"),
	(b"01000010001001110001001100001100", b"01000010101100010111110101101100"), -- 46.9764 + 41.7686 = 88.745
	(b"11000010101001100111101101001100", b"00000000000000000000000000000000"),
	(b"01000001101101011001001001111100", b"11000010011100100010110101011010"), -- -83.2408 + 22.6965 = -60.5443
	(b"10111111111100000111111000000000", b"00000000000000000000000000000000"),
	(b"11000010110000101010000100000100", b"11000010110001100110001011111100"), -- -1.87885 + -97.3145 = -99.1933
	(b"11000010011111110111100001011100", b"00000000000000000000000000000000"),
	(b"01000000101011110001101011100000", b"11000010011010011001010100000000"), -- -63.8675 + 5.47203 = -58.3955
	(b"11000010000110110111111001001011", b"00000000000000000000000000000000"),
	(b"01000001110000001100111111000100", b"11000001011011000101100110100100"), -- -38.8733 + 24.1014 = -14.7719
	(b"11000010001111011110111000010000", b"00000000000000000000000000000000"),
	(b"01000010101011100011011100010000", b"01000010000111101000000000010000"), -- -47.4825 + 87.1075 = 39.6251
	(b"11000010101100010100100100100101", b"00000000000000000000000000000000"),
	(b"01000010101000011110011101000011", b"11000000111101100001111000100000"), -- -88.6429 + 80.9517 = -7.69118
	(b"01000010101110111111001000001000", b"00000000000000000000000000000000"),
	(b"11000010000010011000010111111000", b"01000010011011100101111000011000"), -- 93.9727 + -34.3808 = 59.5919
	(b"01000010100010111110110101111110", b"00000000000000000000000000000000"),
	(b"11000010100101110111100111110100", b"11000000101110001100011101100000"), -- 69.9639 + -75.7382 = -5.77434
	(b"01000010101001110100000000101100", b"00000000000000000000000000000000"),
	(b"11000001010001010110111010101000", b"01000010100011101001001001010111"), -- 83.6253 + -12.3395 = 71.2858
	(b"11000010000101100010001110100100", b"00000000000000000000000000000000"),
	(b"11000010100100011011001111111000", b"11000010110111001100010111001010"), -- -37.5348 + -72.8515 = -110.386
	(b"11000001101001011101111110011100", b"00000000000000000000000000000000"),
	(b"01000010011001000110010110011100", b"01000010000100010111010111001110"), -- -20.7342 + 57.0992 = 36.365
	(b"11000000111001011110110111000000", b"00000000000000000000000000000000"),
	(b"11000010100011010011000000111110", b"11000010100110111000111100011010"), -- -7.18527 + -70.5942 = -77.7795
	(b"11000010101011000011111011100100", b"00000000000000000000000000000000"),
	(b"11000010001000111100000010110111", b"11000010111111100001111101000000"), -- -86.1228 + -40.9382 = -127.061
	(b"11000001100010101010010010001100", b"00000000000000000000000000000000"),
	(b"01000010100001110001101101101100", b"01000010010010001110010010010010"), -- -17.3303 + 67.5536 = 50.2232
	(b"11000010001101111001011010110100", b"00000000000000000000000000000000"),
	(b"01000010110000110011111111111000", b"01000010010011101110100100111100"), -- -45.8972 + 97.6249 = 51.7278
	(b"01000010000110010101111001111100", b"00000000000000000000000000000000"),
	(b"01000001111111101000000111101100", b"01000010100011000100111110111001"), -- 38.3423 + 31.8134 = 70.1557
	(b"01000001111001101111000101101000", b"00000000000000000000000000000000"),
	(b"11000010100100001001100100100010", b"11000010001011011011100110010000"), -- 28.8679 + -72.2991 = -43.4312
	(b"11000010100011001110111001000111", b"00000000000000000000000000000000"),
	(b"11000010011011011001101100110100", b"11000011000000011101110111110000"), -- -70.4654 + -59.4016 = -129.867
	(b"01000001000110110100101101100000", b"00000000000000000000000000000000"),
	(b"11000010100000010111111001101110", b"11000010010111000010101000000100"), -- 9.7059 + -64.7469 = -55.041
	(b"11000010100010110010010101000100", b"00000000000000000000000000000000"),
	(b"11000010100101111101110001101010", b"11000011000100011000000011010111"), -- -69.5728 + -75.9305 = -145.503
	(b"11000001100010111100101011100100", b"00000000000000000000000000000000"),
	(b"11000000101010010010100000000000", b"11000001101101100001010011100100"), -- -17.4741 + -5.28613 = -22.7602
	(b"11000010001011110111001111100000", b"00000000000000000000000000000000"),
	(b"11000010101010001001110100011100", b"11000011000000000010101110000110"), -- -43.8632 + -84.3069 = -128.17
	(b"01000001100001100000011101000000", b"00000000000000000000000000000000"),
	(b"01000010101011001101110001101110", b"01000010110011100101111000111110"), -- 16.7535 + 86.4305 = 103.184
	(b"11000010011111101000001100001000", b"00000000000000000000000000000000"),
	(b"01000010101111111111111000110111", b"01000010000000010111100101100110"), -- -63.628 + 95.9965 = 32.3686
	(b"11000000100000010110000110000000", b"00000000000000000000000000000000"),
	(b"11000010101011111011110010010000", b"11000010101101111101001010101000"), -- -4.04315 + -87.8683 = -91.9114
	(b"01000010010110000001000111101010", b"00000000000000000000000000000000"),
	(b"01000010001110000110011101000110", b"01000010110010000011110010011000"), -- 54.0175 + 46.1009 = 100.118
	(b"01000000101101100100110011100000", b"00000000000000000000000000000000"),
	(b"01000010011000001000001011111110", b"01000010011101110100110010011010"), -- 5.69688 + 56.1279 = 61.8248
	(b"01000010000110111111001001011100", b"00000000000000000000000000000000"),
	(b"11000010100100100111100011101000", b"11000010000010001111111101110100"), -- 38.9867 + -73.2361 = -34.2495
	(b"11000010100110101010100100011000", b"00000000000000000000000000000000"),
	(b"11000010011000101110010011000101", b"11000011000001100000110110111101"), -- -77.3303 + -56.7234 = -134.054
	(b"11000010001111000110110100110000", b"00000000000000000000000000000000"),
	(b"11000001111011010101101111111000", b"11000010100110011000110110010110"), -- -47.1066 + -29.6699 = -76.7765
	(b"01000010000011110100110100011110", b"00000000000000000000000000000000"),
	(b"11000010110001001001111111101100", b"11000010011110011111001010111010"), -- 35.8253 + -98.3123 = -62.487
	(b"01000001110010101000110010010000", b"00000000000000000000000000000000"),
	(b"10111111011000100010001110000000", b"01000001110000110111101101110100"), -- 25.3186 + -0.883354 = 24.4353
	(b"11000010100010100000110000101110", b"00000000000000000000000000000000"),
	(b"11000001110001010011101000111100", b"11000010101110110101101010111101"), -- -69.0238 + -24.6534 = -93.6772
	(b"11000001101001110011110111111100", b"00000000000000000000000000000000"),
	(b"01000001110011100011010011100000", b"01000000100110111101101110010000"), -- -20.9053 + 25.7758 = 4.87055
	(b"11000010000010100000100001011000", b"00000000000000000000000000000000"),
	(b"00111111110001110110001000000000", b"11000010000000111100110101001000"), -- -34.5081 + 1.55768 = -32.9505
	(b"01000010010100100000001011101000", b"00000000000000000000000000000000"),
	(b"11000001000011100001001010110000", b"01000010001011100111111000111100"), -- 52.5028 + -8.87956 = 43.6233
	(b"01000010100100000011011110100111", b"00000000000000000000000000000000"),
	(b"11000001011000010111100100110000", b"01000010011010000001000100000010"), -- 72.1087 + -14.0921 = 58.0166
	(b"01000010001101101000000011111010", b"00000000000000000000000000000000"),
	(b"01000010100101001111010000010110", b"01000010111100000011010010010011"), -- 45.626 + 74.4767 = 120.103
	(b"11000010001111011010000000010110", b"00000000000000000000000000000000"),
	(b"01000001000000010110110111000000", b"11000010000111010100010010100110"), -- -47.4063 + 8.08929 = -39.317
	(b"01000010101001100001100101011111", b"00000000000000000000000000000000"),
	(b"11000010100001111010000000001100", b"01000001011100111100101010011000"), -- 83.0496 + -67.8126 = 15.237
	(b"11000001011000110100011110001000", b"00000000000000000000000000000000"),
	(b"11000010100000011010110100100100", b"11000010100111100001011000010101"), -- -14.205 + -64.8382 = -79.0431
	(b"01000010001010000100110111010010", b"00000000000000000000000000000000"),
	(b"01000010100000110001101011011010", b"01000010110101110100000111000011"), -- 42.076 + 65.5524 = 107.628
	(b"11000010010011000100001000101101", b"00000000000000000000000000000000"),
	(b"01000010101110000011001100101010", b"01000010001001000010010000100111"), -- -51.0646 + 92.0999 = 41.0353
	(b"01000010101000001001100001100101", b"00000000000000000000000000000000"),
	(b"11000001011000101010010101010000", b"01000010100001000100001110111011"), -- 80.2976 + -14.1654 = 66.1323
	(b"01000010110000100000010101011111", b"00000000000000000000000000000000"),
	(b"01000010101001001001011010000010", b"01000011001100110100110111110000"), -- 97.0105 + 82.294 = 179.304
	(b"11000010100010111111011001111100", b"00000000000000000000000000000000"),
	(b"11000001001101000100111000010000", b"11000010101000101000000000111110"), -- -69.9814 + -11.2691 = -81.2505
	(b"01000000010111100101101001100000", b"00000000000000000000000000000000"),
	(b"01000001101001100111001011101000", b"01000001110000100011111000110100"), -- 3.47427 + 20.8061 = 24.2804
	(b"01000010001111001101000110100100", b"00000000000000000000000000000000"),
	(b"01000010110000110100000011111000", b"01000011000100001101010011100101"), -- 47.2047 + 97.6269 = 144.832
	(b"01000010100010110011010101001010", b"00000000000000000000000000000000"),
	(b"11000010101100101100101000110011", b"11000001100111100101001110100100"), -- 69.6041 + -89.3949 = -19.7908
	(b"01000001100110001101100011101000", b"00000000000000000000000000000000"),
	(b"01000010101011001110010111100010", b"01000010110100110001110000011100"), -- 19.1059 + 86.449 = 105.555
	(b"01000001000110001010011110100000", b"00000000000000000000000000000000"),
	(b"11000010000111100100011101000110", b"11000001111100000011101010111100"), -- 9.54092 + -39.5696 = -30.0287
	(b"01000001110000011100111100101000", b"00000000000000000000000000000000"),
	(b"01000001100010101111011011000000", b"01000010001001100110001011110100"), -- 24.2262 + 17.3705 = 41.5966
	(b"11000001110101000010101000000000", b"00000000000000000000000000000000"),
	(b"01000001101100001011010110011100", b"11000000100011011101000110010000"), -- -26.5205 + 22.0887 = -4.43183
	(b"01000010010011100001000101101000", b"00000000000000000000000000000000"),
	(b"11000001001111101001000001110000", b"01000010000111100110110101001100"), -- 51.517 + -11.9103 = 39.6067
	(b"01000001101011000101010100101000", b"00000000000000000000000000000000"),
	(b"11000010101111101000111010000110", b"11000010100100110111100100111100"), -- 21.5416 + -95.2784 = -73.7368
	(b"01000010011001011001000000101101", b"00000000000000000000000000000000"),
	(b"01000010101110101000001101001100", b"01000011000101101010010110110001"), -- 57.3908 + 93.2564 = 150.647
	(b"11000010010100110001111001100110", b"00000000000000000000000000000000"),
	(b"01000010000110111110100110011000", b"11000001010111001101001100111000"), -- -52.7797 + 38.9781 = -13.8016
	(b"11000010110001111111010101100110", b"00000000000000000000000000000000"),
	(b"11000010001011110110011011111110", b"11000011000011111101010001110010"), -- -99.9793 + -43.8506 = -143.83
	(b"11000010100001011101000111101011", b"00000000000000000000000000000000"),
	(b"01000010110001011101111111010011", b"01000010000000000001101111010000"), -- -66.91 + 98.9372 = 32.0272
	(b"01000010100011000110000101101100", b"00000000000000000000000000000000"),
	(b"11000001010101100111000010000000", b"01000010011000110010011010111000"), -- 70.1903 + -13.4025 = 56.7878
	(b"11000010000010010100011100010100", b"00000000000000000000000000000000"),
	(b"01000010001010011011001001010110", b"01000001000000011010110100001000"), -- -34.3194 + 42.4242 = 8.10474
	(b"01000010101011010111101010110010", b"00000000000000000000000000000000"),
	(b"01000001110100000101011001110100", b"01000010111000011001000001001111"), -- 86.7396 + 26.0422 = 112.782
	(b"01000010100001111101100110000010", b"00000000000000000000000000000000"),
	(b"11000000011111101001011010100000", b"01000010011111111100100110011010"), -- 67.9248 + -3.97794 = 63.9469
	(b"11000001000011001111111100111000", b"00000000000000000000000000000000"),
	(b"01000001101101001101001110001000", b"01000001010111001010011111011000"), -- -8.81231 + 22.6033 = 13.791
	(b"01000001100000000101010111000100", b"00000000000000000000000000000000"),
	(b"01000010100001010111111101010110", b"01000010101001011001010011000111"), -- 16.0419 + 66.7487 = 82.7906
	(b"11000010100001111111110101110100", b"00000000000000000000000000000000"),
	(b"01000010101000110001000110111110", b"01000001010110001010001001010000"), -- -67.995 + 81.5347 = 13.5396
	(b"01000010010010010000011110110100", b"00000000000000000000000000000000"),
	(b"11000000110000001110100010110000", b"01000010001100001110101010011110"), -- 50.2575 + -6.0284 = 44.2291
	(b"11000000111000101100100000110000", b"00000000000000000000000000000000"),
	(b"11000010100001111111111010101010", b"11000010100101100010101100101101"), -- -7.08694 + -67.9974 = -75.0843
	(b"01000001000010101001101110000000", b"00000000000000000000000000000000"),
	(b"11000001101000000111101000000000", b"11000001001101100101100010000000"), -- 8.66296 + -20.0596 = -11.3966
	(b"11000010101001010110010110111000", b"00000000000000000000000000000000"),
	(b"11000001110100110100111101010000", b"11000010110110100011100110001100"), -- -82.6987 + -26.4137 = -109.112
	(b"11000010101101000110001110010010", b"00000000000000000000000000000000"),
	(b"01000001101010010110110000111000", b"11000010100010100000100010000100"), -- -90.1945 + 21.1778 = -69.0166
	(b"01000010100000010010000010011100", b"00000000000000000000000000000000"),
	(b"11000001101000011100000111011100", b"01000010001100010110000001001010"), -- 64.5637 + -20.2197 = 44.344
	(b"11000010101100000011010011100100", b"00000000000000000000000000000000"),
	(b"11000000111110101100111100110000", b"11000010101111111110000111010111"), -- -88.1033 + -7.83779 = -95.9411
	(b"11000010000001011000001011111100", b"00000000000000000000000000000000"),
	(b"01000010101010110111100011001010", b"01000010010100010110111010011000"), -- -33.3779 + 85.7359 = 52.358
	(b"01000010100011110110101001100010", b"00000000000000000000000000000000"),
	(b"01000010101111010001100110001000", b"01000011001001100100000111110101"), -- 71.7078 + 94.5499 = 166.258
	(b"01000010101000010011001001111101", b"00000000000000000000000000000000"),
	(b"01000010001100000110110011010000", b"01000010111110010110100011100101"), -- 80.5986 + 44.1063 = 124.705
	(b"11000010101110000000100000010101", b"00000000000000000000000000000000"),
	(b"01000010100010110000111110011110", b"11000001101100111110000111011100"), -- -92.0158 + 69.5305 = -22.4853
	(b"11000000111000010110100101100000", b"00000000000000000000000000000000"),
	(b"11000001000100010011010110010000", b"11000001100000001111010100100000"), -- -7.04411 + -9.07558 = -16.1197
	(b"01000001101011110011010111011000", b"00000000000000000000000000000000"),
	(b"11000001110000110011100010001100", b"11000000001000000001010110100000"), -- 21.9013 + -24.4026 = -2.50132
	(b"11000010100100101110000001110110", b"00000000000000000000000000000000"),
	(b"01000000010011010110111110100000", b"11000010100011000111010011111001"), -- -73.4384 + 3.20994 = -70.2285
	(b"01000010010111010111010101000100", b"00000000000000000000000000000000"),
	(b"11000010011001010000101100111000", b"10111111111100101011111010000000"), -- 55.3645 + -57.261 = -1.89644
	(b"11000010100010101100110110111001", b"00000000000000000000000000000000"),
	(b"11000010100100100110011100110110", b"11000011000011101001101001111000"), -- -69.4018 + -73.2016 = -142.603
	(b"11000001010110010100011010011000", b"00000000000000000000000000000000"),
	(b"01000001011111111001011011100000", b"01000000000110010100000100100000"), -- -13.5797 + 15.9743 = 2.3946
	(b"01000010101001010000011111010110", b"00000000000000000000000000000000"),
	(b"01000010011110000011110111110100", b"01000011000100001001001101101000"), -- 82.5153 + 62.0605 = 144.576
	(b"01000010100001110110100101101010", b"00000000000000000000000000000000"),
	(b"01000010100110011110011001001000", b"01000011000100001010011111011001"), -- 67.7059 + 76.9498 = 144.656
	(b"11000010010100001100011010011010", b"00000000000000000000000000000000"),
	(b"11000010101100110110001000010010", b"11000011000011011110001010110000"), -- -52.1939 + -89.6915 = -141.885
	(b"01000010101111000010010100101110", b"00000000000000000000000000000000"),
	(b"11000010100100011101000110101100", b"01000001101010010100111000001000"), -- 94.0726 + -72.9095 = 21.1631
	(b"01000010001011010101100010011000", b"00000000000000000000000000000000"),
	(b"11000010101111001110000101010010", b"11000010010011000110101000001100"), -- 43.3365 + -94.4401 = -51.1036
	(b"11000001000101111011100110101000", b"00000000000000000000000000000000"),
	(b"11000010010011001000101111111000", b"11000010011100100111101001100010"), -- -9.48283 + -51.1367 = -60.6195
	(b"11000000011110110101100000100000", b"00000000000000000000000000000000"),
	(b"01000010101010101011101000011000", b"01000010101000101101111101010111"), -- -3.92725 + 85.3635 = 81.4362
	(b"01000010011010110101000110000011", b"00000000000000000000000000000000"),
	(b"01000001011010010101101000111000", b"01000010100100101101010000001000"), -- 58.8296 + 14.5845 = 73.4141
	(b"11000010100111101001101010000110", b"00000000000000000000000000000000"),
	(b"11000001101101110011110110111100", b"11000010110011000110100111110101"), -- -79.3018 + -22.9051 = -102.207
	(b"01000010000110101000111101001100", b"00000000000000000000000000000000"),
	(b"01000010011010111100110010100000", b"01000010110000110010110111110110"), -- 38.6399 + 58.9498 = 97.5898
	(b"01000010010010001100001011000000", b"00000000000000000000000000000000"),
	(b"11000010110000010000010011001000", b"11000010001110010100011011010000"), -- 50.1902 + -96.5093 = -46.3192
	(b"10111110011101111100000000000000", b"00000000000000000000000000000000"),
	(b"11000001100011100000110001000000", b"11000001100011111111101111000000"), -- -0.241943 + -17.756 = -17.9979
	(b"11000010101111011111001010000110", b"00000000000000000000000000000000"),
	(b"11000001001110011101010011001000", b"11000010110101010010110100011111"), -- -94.9737 + -11.6144 = -106.588
	(b"11000010011100001111110100110011", b"00000000000000000000000000000000"),
	(b"01000001100010101010011101100100", b"11000010001010111010100110000001"), -- -60.2473 + 17.3317 = -42.9155
	(b"11000001111100110111010111111000", b"00000000000000000000000000000000"),
	(b"11000010100110110111011100000011", b"11000010110110000101010010000001"), -- -30.4326 + -77.7324 = -108.165
	(b"01000001110001011011110100100000", b"00000000000000000000000000000000"),
	(b"11000001101000101110111111011000", b"01000000100010110011010100100000"), -- 24.7173 + -20.3671 = 4.35023
	(b"01000010100010001010101001010110", b"00000000000000000000000000000000"),
	(b"01000010101000110000000100101010", b"01000011000101011101010111000000"), -- 68.3327 + 81.5023 = 149.835
	(b"01000010000010111011111000011010", b"00000000000000000000000000000000"),
	(b"01000010100111100001001000110011", b"01000010111000111111000101000000"), -- 34.9356 + 79.0355 = 113.971
	(b"01000001110001100100000000101100", b"00000000000000000000000000000000"),
	(b"01000001111111010110101000100100", b"01000010011000011101010100101000"), -- 24.7813 + 31.6768 = 56.4582
	(b"01000010110001001000100011100000", b"00000000000000000000000000000000"),
	(b"01000010010100000011111001001110", b"01000011000101100101010000000100"), -- 98.2673 + 52.0608 = 150.328
	(b"11000010101011001000100011100001", b"00000000000000000000000000000000"),
	(b"01000010101011011010000010100000", b"00111111000010111101111110000000"), -- -86.2673 + 86.8137 = 0.546379
	(b"11000001111111010100011100000000", b"00000000000000000000000000000000"),
	(b"01000010010001010001001001101000", b"01000001100011001101110111010000"), -- -31.6597 + 49.268 = 17.6083
	(b"01000010001100100000110110010100", b"00000000000000000000000000000000"),
	(b"11000000000100010111100000000000", b"01000010001010001111011000010100"), -- 44.5133 + -2.27295 = 42.2403
	(b"11000000011000010001110100000000", b"00000000000000000000000000000000"),
	(b"11000010100001000110010101111010", b"11000010100010110110111001100010"), -- -3.5174 + -66.1982 = -69.7156
	(b"01000010001011001011010011010000", b"00000000000000000000000000000000"),
	(b"11000000010011101010111010000000", b"01000010000111111100100111101000"), -- 43.1766 + -3.2294 = 39.9472
	(b"01000010011111000010000101111100", b"00000000000000000000000000000000"),
	(b"01000001101111111101101110011000", b"01000010101011100000011110100100"), -- 63.0327 + 23.9822 = 87.0149
	(b"11000010011110001011101000101101", b"00000000000000000000000000000000"),
	(b"01000010010010010101000000100111", b"11000001001111011010100000011000"), -- -62.1818 + 50.3283 = -11.8535
	(b"01000001110111011101010111001100", b"00000000000000000000000000000000"),
	(b"01000010101011111011001011110000", b"01000010111001110010100001100011"), -- 27.7294 + 87.8495 = 115.579
	(b"11000001101101010111101100101000", b"00000000000000000000000000000000"),
	(b"11000010001010011110011111010100", b"11000010100000100101001010110100"), -- -22.6851 + -42.4764 = -65.1615
	(b"11000010100000111000001100100000", b"00000000000000000000000000000000"),
	(b"11000010011100010000001100101101", b"11000010111111000000010010110110"), -- -65.7561 + -60.2531 = -126.009
	(b"01000001100011011000111011010000", b"00000000000000000000000000000000"),
	(b"11000010011111011011101111010111", b"11000010001101101111010001101111"), -- 17.6947 + -63.4334 = -45.7387
	(b"11000010101100100100000010100000", b"00000000000000000000000000000000"),
	(b"11000001011000011010001000111000", b"11000010110011100111010011100111"), -- -89.1262 + -14.1021 = -103.228
	(b"01000010011010110100111010111000", b"00000000000000000000000000000000"),
	(b"11000001001011000000100010010000", b"01000010010000000100110010010100"), -- 58.8269 + -10.7521 = 48.0748
	(b"01000010101010001110011100100010", b"00000000000000000000000000000000"),
	(b"11000001110101111111100111100000", b"01000010011001011101000101010100"), -- 84.4514 + -26.997 = 57.4544
	(b"01000010011110111010101010101010", b"00000000000000000000000000000000"),
	(b"11000010101101011101110010100000", b"11000001111000000001110100101100"), -- 62.9167 + -90.9309 = -28.0142
	(b"01000001110111001001011011111000", b"00000000000000000000000000000000"),
	(b"11000010001101111000101010010111", b"11000001100100100111111000110110"), -- 27.5737 + -45.8853 = -18.3116
	(b"01000010100110111011000011000110", b"00000000000000000000000000000000"),
	(b"11000001110101110111010000100000", b"01000010010010111010011101111100"), -- 77.8453 + -26.9317 = 50.9136
	(b"11000001000011100001101101010000", b"00000000000000000000000000000000"),
	(b"11000010011100101001011101111000", b"11000010100010110000111100100110"), -- -8.88167 + -60.6479 = -69.5296
	(b"01000001110001000011011011010100", b"00000000000000000000000000000000"),
	(b"11000010000000000100001111101010", b"11000000111100010100010000000000"), -- 24.5268 + -32.0663 = -7.53955
	(b"11000010001111101111000101010100", b"00000000000000000000000000000000"),
	(b"01000010100101000000111001111100", b"01000001110100100101011101001000"), -- -47.7357 + 74.0283 = 26.2926
	(b"11000010100101111110101000011000", b"00000000000000000000000000000000"),
	(b"11000010100101010111011000011111", b"11000011000101101011000000011100"), -- -75.9572 + -74.7307 = -150.688
	(b"01000010100100100100100001101011", b"00000000000000000000000000000000"),
	(b"01000001010100010010010100000000", b"01000010101011000110110100001011"), -- 73.1414 + 13.0715 = 86.213
	(b"11000010110000110101010110011000", b"00000000000000000000000000000000"),
	(b"01000010000100000000000111100000", b"11000010011101101010100101010000"), -- -97.6672 + 36.0018 = -61.6653
	(b"01000010100100010111011000110000", b"00000000000000000000000000000000"),
	(b"11000010010101011110100100101000", b"01000001100110100000011001110000"), -- 72.7308 + -53.4777 = 19.2531
	(b"01000010100010010000111000010010", b"00000000000000000000000000000000"),
	(b"11000001001101101111110110011000", b"01000010011001000101110010111110"), -- 68.5275 + -11.4369 = 57.0906
	(b"01000010001000010100001101011010", b"00000000000000000000000000000000"),
	(b"01000010011100110110000011100001", b"01000010110010100101001000011110"), -- 40.3158 + 60.8446 = 101.16
	(b"01000001010010111011100001110000", b"00000000000000000000000000000000"),
	(b"11000010100010100100110111110000", b"11000010011000011010110111000100"), -- 12.7325 + -69.1522 = -56.4197
	(b"11000000101011001000111111100000", b"00000000000000000000000000000000"),
	(b"01000010011000101101101001101000", b"01000010010011010100100001101100"), -- -5.39256 + 56.7133 = 51.3207
	(b"01000010001100111001010001000110", b"00000000000000000000000000000000"),
	(b"11000001101001101111101011110100", b"01000001110000000010110110011000"), -- 44.8948 + -20.8725 = 24.0223
	(b"01000010010011110011001011000111", b"00000000000000000000000000000000"),
	(b"01000010101001011100001101101001", b"01000011000001101010111001100110"), -- 51.7996 + 82.8817 = 134.681
	(b"01000010001100110110111010101110", b"00000000000000000000000000000000"),
	(b"11000010101010001101101001101100", b"11000010000111100100011000101010"), -- 44.8581 + -84.4266 = -39.5685
	(b"11000000111110111011111010010000", b"00000000000000000000000000000000"),
	(b"11000001111001001010001100001000", b"11000010000100011100100101010110"), -- -7.86701 + -28.5796 = -36.4466
	(b"01000010100011010010101100010100", b"00000000000000000000000000000000"),
	(b"01000000011011110101000101100000", b"01000010100101001010010110011111"), -- 70.5841 + 3.73934 = 74.3235
	(b"01000001100011010110110001001000", b"00000000000000000000000000000000"),
	(b"01000001110011111111010011000100", b"01000010001011101011000010000110"), -- 17.6779 + 25.9945 = 43.6724
	(b"01000000001101001101111000000000", b"00000000000000000000000000000000"),
	(b"11000001101101100001111010010100", b"11000001100111111000001011010100"), -- 2.82605 + -22.7649 = -19.9389
	(b"01000010100101100011011101011101", b"00000000000000000000000000000000"),
	(b"01000010100011111110001010111000", b"01000011000100110000110100001010"), -- 75.1081 + 71.9428 = 147.051
	(b"10111101110000110110010000000000", b"00000000000000000000000000000000"),
	(b"01000001000110010100000101011000", b"01000001000101111011101010010000"), -- -0.0954056 + 9.57845 = 9.48305
	(b"01000001001100110001101011100000", b"00000000000000000000000000000000"),
	(b"01000010100101101110110001001010", b"01000010101011010100111110100110"), -- 11.1941 + 75.4615 = 86.6556
	(b"01000010010000110110100111110101", b"00000000000000000000000000000000"),
	(b"01000010011011000101000011011000", b"01000010110101111101110101100110"), -- 48.8535 + 59.0789 = 107.932
	(b"11000010100011000111001000011100", b"00000000000000000000000000000000"),
	(b"11000001110010100111110010100100", b"11000010101111110001000101000101"), -- -70.2229 + -25.3109 = -95.5337
	(b"11000010100111000001011010100100", b"00000000000000000000000000000000"),
	(b"11000010011010001000011100101000", b"11000011000010000010110100011100"), -- -78.0442 + -58.132 = -136.176
	(b"01000010001110101000000010101100", b"00000000000000000000000000000000"),
	(b"11000010011011111111100101001100", b"11000001010101011110001010000000"), -- 46.6257 + -59.9935 = -13.3678
	(b"01000001110010000001111101111000", b"00000000000000000000000000000000"),
	(b"01000010011010100111100010010100", b"01000010101001110100010000101000"), -- 25.0154 + 58.6178 = 83.6331
	(b"11000010001010000011110000000000", b"00000000000000000000000000000000"),
	(b"01000001110110010111011011110000", b"11000001011011100000001000100000"), -- -42.0586 + 27.1831 = -14.8755
	(b"01000001100011011100110111010000", b"00000000000000000000000000000000"),
	(b"01000010011111101100111011010100", b"01000010101000101101101011011110"), -- 17.7255 + 63.702 = 81.4275
	(b"11000001010000100011101001000000", b"00000000000000000000000000000000"),
	(b"01000010101011001000110011100001", b"01000010100101000100010110011001"), -- -12.1392 + 86.2752 = 74.1359
	(b"11000010101101111111010110010010", b"00000000000000000000000000000000"),
	(b"00111110011001101101100000000000", b"11000010101101111000001000100110"), -- -91.9796 + 0.225433 = -91.7542
	(b"01000001101000011100000000000100", b"00000000000000000000000000000000"),
	(b"11000000101000010010010110110000", b"01000001011100101110110100110000"), -- 20.2188 + -5.03585 = 15.1829
	(b"11000001110101101101000101101000", b"00000000000000000000000000000000"),
	(b"11000010001101011001110111001011", b"11000010100100001000001101000000"), -- -26.8522 + -45.4041 = -72.2563
	(b"01000010101101001101001000000010", b"00000000000000000000000000000000"),
	(b"01000010101100000001010111101000", b"01000011001100100111001111110101"), -- 90.4102 + 88.0428 = 178.453
	(b"10110100000000011010110010101011", b"00000000000000000000000000000000"),
	(b"11000010011010111011110111111100", b"11000010011010111011110111111100"), -- -1.20769e-07 + -58.9355 = -58.9355
	(b"10011010111010000110000110110000", b"00000000000000000000000000000000"),
	(b"10110111100100010010000110010010", b"10110111100100010010000110010010"), -- -9.61108e-23 + -1.7301e-05 = -1.7301e-05
	(b"11000010101000100110001010011111", b"00000000000000000000000000000000"),
	(b"10110111101100001101000011100010", b"11000010101000100110001010100010"), -- -81.1926 + -2.10781e-05 = -81.1926
	(b"10101001000010110101001100110100", b"00000000000000000000000000000000"),
	(b"11000110001011000001110101111011", b"11000110001011000001110101111011"), -- -3.09364e-14 + -11015.4 = -11015.4
	(b"01001010001000100101011111000011", b"00000000000000000000000000000000"),
	(b"10101111111001110001110101010011", b"01001010001000100101011111000011"), -- 2.65982e+06 + -4.20395e-10 = 2.65982e+06
	(b"00111010101001011011000010000010", b"00000000000000000000000000000000"),
	(b"00111110110111011010100110111000", b"00111110110111100100111101101001"), -- 0.00126411 + 0.432935 = 0.4342
	(b"10110101100010100101010000010011", b"00000000000000000000000000000000"),
	(b"11001111110011111101101100101000", b"11001111110011111101101100101000"), -- -1.03063e-06 + -6.97449e+09 = -6.97449e+09
	(b"11000101001000101100011001000000", b"00000000000000000000000000000000"),
	(b"01001010010100111110011101000111", b"01001010010100111011111010010101"), -- -2604.39 + 3.47183e+06 = 3.46922e+06
	(b"01001100110001110100001010101001", b"00000000000000000000000000000000"),
	(b"01010011001000110011010110011000", b"01010011001000110011101111010010"), -- 1.0447e+08 + 7.00979e+11 = 7.01083e+11
	(b"11000000011111101110010010101011", b"00000000000000000000000000000000"),
	(b"11010100000111000010101101111101", b"11010100000111000010101101111101"), -- -3.98271 + -2.68298e+12 = -2.68298e+12
	(b"00110000010101000101101110100101", b"00000000000000000000000000000000"),
	(b"10101010000000000000000100100011", b"00110000010101000101001110100101"), -- 7.72554e-10 + -1.13691e-13 = 7.7244e-10
	(b"00111100001100000110000001000101", b"00000000000000000000000000000000"),
	(b"10110101101110100110011100001101", b"00111100001100000101101001110010"), -- 0.0107651 + -1.38881e-06 = 0.0107638
	(b"00111100101001011011111001100110", b"00000000000000000000000000000000"),
	(b"11010101011000101001111011111000", b"11010101011000101001111011111000"), -- 0.0202324 + -1.55733e+13 = -1.55733e+13
	(b"11000101010101011010001110010001", b"00000000000000000000000000000000"),
	(b"00110010001000011001100110000011", b"11000101010101011010001110010001"), -- -3418.22 + 9.40634e-09 = -3418.22
	(b"10010001110000000010101111101111", b"00000000000000000000000000000000"),
	(b"01000101100101101100101100111000", b"01000101100101101100101100111000"), -- -3.03193e-28 + 4825.4 = 4825.4
	(b"00111010011100111011111111110100", b"00000000000000000000000000000000"),
	(b"00101110000111100010011100000111", b"00111010011100111011111111110101"), -- 0.000929832 + 3.59597e-11 = 0.000929832
	(b"01001100101111110101101111101111", b"00000000000000000000000000000000"),
	(b"11000111001010110110001001001101", b"01001100101111110100011010000011"), -- 1.00327e+08 + -43874.3 = 1.00283e+08
	(b"00100101101001000101101010110011", b"00000000000000000000000000000000"),
	(b"01010010000100100101110110101101", b"01010010000100100101110110101101"), -- 2.85109e-16 + 1.57159e+11 = 1.57159e+11
	(b"11010110100100000101001111011100", b"00000000000000000000000000000000"),
	(b"11010010100110101100110011111100", b"11010110100100001110111010101001"), -- -7.93449e+13 + -3.32432e+11 = -7.96774e+13
	(b"11000000001101010001001111001111", b"00000000000000000000000000000000"),
	(b"10110000100011100000000111100000", b"11000000001101010001001111001111"), -- -2.82933 + -1.03324e-09 = -2.82933
	(b"00110000001011011100100100001001", b"00000000000000000000000000000000"),
	(b"00111010111010001011110110001111", b"00111010111010001011110110010100"), -- 6.32227e-10 + 0.00177567 = 0.00177567
	(b"01000010010000010000110011100101", b"00000000000000000000000000000000"),
	(b"00111000110010010100111010101111", b"01000010010000010000110011111110"), -- 48.2626 + 9.59908e-05 = 48.2627
	(b"11001101110000001111111110011110", b"00000000000000000000000000000000"),
	(b"10101001000010111001110100011000", b"11001101110000001111111110011110"), -- -4.04747e+08 + -3.10005e-14 = -4.04747e+08
	(b"11011001001101101111111111111111", b"00000000000000000000000000000000"),
	(b"10110010101000011000100011100011", b"11011001001101101111111111111111"), -- -3.21937e+15 + -1.88051e-08 = -3.21937e+15
	(b"00111111111011011011010110111000", b"00000000000000000000000000000000"),
	(b"01000001001101111000110111010011", b"01000001010101010100010010001010"), -- 1.85711 + 11.4721 = 13.3292
	(b"11001101011111010000001000110001", b"00000000000000000000000000000000"),
	(b"11001110110101001001111000001011", b"11001110111101000011111001010001"), -- -2.65299e+08+-1.78356e+09=-2.04886e+09
	(b"01001100111011111110101010101111", b"00000000000000000000000000000000"),
	(b"11001110101110001101010010001101", b"11001110101010011101010111100010"), -- 1.25785e+08+-1.55047e+09=-1.42468e+09
	(b"11001110100100010110111000100110", b"00000000000000000000000000000000"),
	(b"01001110100010110001001000010111", b"11001100010010111000000111100000"), -- -1.21996e+09+1.16661e+09=-5.33482e+07
	(b"01001110011011011110011010111110", b"00000000000000000000000000000000"),
	(b"11001110110001000000000110011000", b"11001110000110100001110001110010"), -- 9.97831e+08+-1.64422e+09=-6.46389e+08
	(b"01001110000001100101100010011011", b"00000000000000000000000000000000"),
	(b"01001101110000100000001111001000", b"01001110011001110101101001111111"), -- 5.63488e+08+4.06878e+08=9.70367e+08
	(b"01001101100000110000001011101101", b"00000000000000000000000000000000"),
	(b"01001110000110111010111001110011", b"01001110010111010010111111101010"), -- 2.74751e+08+6.52975e+08=9.27726e+08
	(b"11001110111000100101011000100110", b"00000000000000000000000000000000"),
	(b"01001101110000101111010101011011", b"11001110101100011001100011001111"), -- -1.89865e+09+4.08857e+08=-1.48979e+09
	(b"01001101101010100001001110001010", b"00000000000000000000000000000000"),
	(b"11001101101100111101101010101010", b"11001011100111000111001000000000"), -- 3.56676e+08+-3.77182e+08=-2.05056e+07
	(b"01001110011101011001101111001000", b"00000000000000000000000000000000"),
	(b"11001110000101001100111010010111", b"01001101110000011001101001100010"), -- 1.03016e+09+-6.24142e+08=4.06015e+08
	(b"11001110011101100100100101000101", b"00000000000000000000000000000000"),
	(b"01001110000110111010111100000001", b"11001101101101010011010010001000"), -- -1.033e+09+6.52984e+08=-3.80015e+08
	(b"11001110000001001111111010010010", b"00000000000000000000000000000000"),
	(b"11001100011010000101010001111110", b"11001110000100111000001111011010"), -- -5.57819e+08+-6.09039e+07=-6.18723e+08
	(b"01001110101100001001011100000101", b"00000000000000000000000000000000"),
	(b"11001110100111111101011010001110", b"01001101000001100000001110111000"), -- 1.48134e+09+-1.34082e+09=1.40524e+08
	(b"11001101100101110000000011100110", b"00000000000000000000000000000000"),
	(b"11001110101010101110101000100100", b"11001110110100001010101001011110"), -- -3.16677e+08+-1.43374e+09=-1.75041e+09
	(b"01001100111111010011111011111111", b"00000000000000000000000000000000"),
	(b"01001110110000001110110010011000", b"01001110110100001100000010001000"), -- 1.32774e+08+1.61837e+09=1.75114e+09
	(b"01001110101110101111000010001001", b"00000000000000000000000000000000"),
	(b"11001110110101001001010111000011", b"11001101010011010010100111010000"), -- 1.56816e+09+-1.78329e+09=-2.15129e+08
	(b"11001011010001100011011011000100", b"00000000000000000000000000000000"),
	(b"11001101001111010001110001010001", b"11001101010010010111111110111101"), -- -1.29901e+07+-1.98297e+08=-2.11287e+08
	(b"11001110010001000001010110101100", b"00000000000000000000000000000000"),
	(b"01001110110001111100001000001101", b"01001110010010110110111001101110"), -- -8.22439e+08+1.67569e+09=8.53253e+08
	(b"01001101000110101010001110111001", b"00000000000000000000000000000000"),
	(b"01001110111000000011101111111011", b"01001110111100111001000001110010"), -- 1.62151e+08+1.88101e+09=2.04316e+09
	(b"01001110111101111101111110000101", b"00000000000000000000000000000000"),
	(b"01001110111101010110110000100110", b"01001111011101101010010111010110"), -- 2.07931e+09+2.05875e+09=4.13806e+09
	(b"11001110101111010010111000110011", b"00000000000000000000000000000000"),
	(b"11001110010101010111001100100001", b"11001111000100111111001111100010"), -- -1.58696e+09+-8.95273e+08=-2.48223e+09
	(b"01001110111111010010011101111111", b"00000000000000000000000000000000"),
	(b"11001110010101001010000100001111", b"01001110100100101101011011111000"), -- 2.12361e+09+-8.91831e+08=1.23178e+09
	(b"01001110111011100001000101011010", b"00000000000000000000000000000000"),
	(b"11001110100011101011111010001011", b"01001110001111101010010110011110"), -- 1.99706e+09+-1.19743e+09=7.99631e+08
	(b"01001110110101101010011000011010", b"00000000000000000000000000000000"),
	(b"01001101111110001001110011010100", b"01001111000010100110011010101000"), -- 1.8006e+09+5.21378e+08=2.32198e+09
	(b"01001110101000011000010111000111", b"00000000000000000000000000000000"),
	(b"01001110110110110001001111101001", b"01001111001111100100110011011000"), -- 1.35495e+09+1.83776e+09=3.19271e+09
	(b"11001101010011101001010011100110", b"00000000000000000000000000000000"),
	(b"11001100011100000100110011001011", b"11001101100001010101010000001100"), -- -2.16617e+08+-6.29932e+07=-2.7961e+08
	(b"01001110111001111011111001100001", b"00000000000000000000000000000000"),
	(b"01001110010100110111101110000001", b"01001111001010001011111000010001"), -- 1.94401e+09+8.87022e+08=2.83103e+09
	(b"11001110001111100101001111001101", b"00000000000000000000000000000000"),
	(b"11001110110100110100001100101110", b"11001111000110010011011010001010"), -- -7.98291e+08+-1.7722e+09=-2.57049e+09
	(b"11001101111101111111001011111100", b"00000000000000000000000000000000"),
	(b"01001110011000010100010000100111", b"01001101110010101001010101010010"), -- -5.19987e+08+9.44835e+08=4.24848e+08
	(b"01001110110110101111001010011011", b"00000000000000000000000000000000"),
	(b"01001101010100000000001110010010", b"01001110111101001111001100001101"), -- 1.83667e+09+2.18118e+08=2.05478e+09
	(b"01001110101010001011111011111101", b"00000000000000000000000000000000"),
	(b"01001110101100110001101111111010", b"01001111001011011110110101111100"), -- 1.41554e+09+1.50248e+09=2.91802e+09
	(b"11001110111100010100001100101111", b"00000000000000000000000000000000"),
	(b"01001101110101101011010000001000", b"11001110101110111001011000101101"), -- -2.02386e+09+4.50265e+08=-1.57359e+09
	(b"11001101000001100000011101010111", b"00000000000000000000000000000000"),
	(b"01001101001001111101001010100010", b"01001100000001110010110100101100"), -- -1.40539e+08+1.75975e+08=3.54357e+07
	(b"11001110011001000000001111001010", b"00000000000000000000000000000000"),
	(b"01001110000011111100101000101100", b"11001101101010000111001100111100"), -- -9.56363e+08+6.03098e+08=-3.53266e+08
	(b"01001110000010110001011100111111", b"00000000000000000000000000000000"),
	(b"01001110110101010110001010100110", b"01001111000011010111011100100011"), -- 5.83389e+08+1.79001e+09=2.3734e+09
	(b"01001110010111100100101001110100", b"00000000000000000000000000000000"),
	(b"01001110011011010010010101111010", b"01001110111001011011011111110111"), -- 9.32355e+08+9.94664e+08=1.92702e+09
	(b"01001110100100111111010000000000", b"00000000000000000000000000000000"),
	(b"11001110001011001100100011001011", b"01001101111101100011111001101010"), -- 1.24112e+09+-7.2471e+08=5.16411e+08
	(b"01001101101000011010101000101101", b"00000000000000000000000000000000"),
	(b"01001110010110101010100001111001", b"01001110100101011011111011001000"), -- 3.39036e+08+9.17119e+08=1.25615e+09
	(b"01001101100101011101110100110010", b"00000000000000000000000000000000"),
	(b"01001110101111001110011100101111", b"01001110111000100101111001111100"), -- 3.14288e+08+1.58463e+09=1.89892e+09
	(b"01001110110010011000110111000101", b"00000000000000000000000000000000"),
	(b"01001110101111010110000101100100", b"01001111010000110111011110010100"), -- 1.69076e+09+1.58864e+09=3.27939e+09
	(b"01001101010100110100011110101000", b"00000000000000000000000000000000"),
	(b"11001110110111001000001110111111", b"11001110110000100001101011001010"), -- 2.21543e+08+-1.84981e+09=-1.62827e+09
	(b"11001101100100011010001101010101", b"00000000000000000000000000000000"),
	(b"01001110110111001001110111101010", b"01001110101110000011010100010101"), -- -3.05425e+08+1.85067e+09=1.54524e+09
	(b"01001110101100100000000010010000", b"00000000000000000000000000000000"),
	(b"11001110101011011010001100110101", b"01001100000010111010101101100000"), -- 1.49319e+09+-1.45658e+09=3.66135e+07
	(b"11001101100100001101011111001000", b"00000000000000000000000000000000"),
	(b"01001110100010100110001001111010", b"01001110010011000101100100010000"), -- -3.03758e+08+1.16085e+09=8.57097e+08
	(b"01001110111000001100011011011111", b"00000000000000000000000000000000"),
	(b"11001110100001000111111001000011", b"01001110001110001001000100111000"), -- 1.88556e+09+-1.11143e+09=7.74131e+08
	(b"01001110111100011101001010000000", b"00000000000000000000000000000000"),
	(b"01001110010010100001110100011111", b"01001111001010110111000010001000"), -- 2.02855e+09+8.47727e+08=2.87628e+09
	(b"01001101100001111101011011111000", b"00000000000000000000000000000000"),
	(b"11001110110001101101100101000101", b"11001110101001001110001110000111"), -- 2.84877e+08+-1.66806e+09=-1.38319e+09
	(b"11001110100001000011101010101010", b"00000000000000000000000000000000"),
	(b"01001110100101010011100010110010", b"01001101000001111111000001000000"), -- -1.10922e+09+1.25176e+09=1.42542e+08
	(b"11001110011000110111100011100011", b"00000000000000000000000000000000"),
	(b"01001110001011001011010101111101", b"11001101010110110000110110011000"), -- -9.54088e+08+7.24394e+08=-2.29694e+08
	(b"01001110100001111110111000001010", b"00000000000000000000000000000000"),
	(b"11001110101010100001110001010010", b"11001101100010001011100100100000"), -- 1.14026e+09+-1.42699e+09=-2.86729e+08
	(b"01001100111100101010111000011100", b"00000000000000000000000000000000"),
	(b"01001110101010001111101101101010", b"01001110101110000010011001001100"), -- 1.27234e+08+1.41752e+09=1.54476e+09
	(b"01001110010111111010100101011111", b"00000000000000000000000000000000"),
	(b"11001101111001000010100111100000", b"01001101110110110010100011011110"), -- 9.38105e+08+-4.78494e+08=4.59611e+08
	(b"01001110110011100100001100101010", b"00000000000000000000000000000000"),
	(b"11001101001000000100100000001110", b"01001110101110100011101000101000"), -- 1.73025e+09+-1.68067e+08=1.56219e+09
	(b"11001110010101001100011110000001", b"00000000000000000000000000000000"),
	(b"01001110101111011100000101110001", b"01001110001001101011101101100001"), -- -8.92461e+08+1.59179e+09=6.99324e+08
	(b"11001011111011100101100010101110", b"00000000000000000000000000000000"),
	(b"01001110110101100011111010011110", b"01001110110100101000010100111011"), -- -3.12405e+07+1.79721e+09=1.76597e+09
	(b"01001110111011010011110010111000", b"00000000000000000000000000000000"),
	(b"01001110100010000111010010100011", b"01001111001110101101100010101110"), -- 1.99009e+09+1.14467e+09=3.13476e+09
	(b"11001110000010100011001000001100", b"00000000000000000000000000000000"),
	(b"11001101011101001110101010010110", b"11001110010001110110110010110010"), -- -5.79634e+08+-2.56813e+08=-8.36447e+08
	(b"11001110001011110100111110010101", b"00000000000000000000000000000000"),
	(b"11001110111001100010110010100100", b"11001111000111101110101000110111"), -- -7.35307e+08+-1.93084e+09=-2.66615e+09
	(b"11001110111110100011010110100110", b"00000000000000000000000000000000"),
	(b"11001101111011101100000000011011", b"11001111000110101111001011010110"), -- -2.09891e+09+-5.00696e+08=-2.59961e+09
	(b"01001110111110010111000101110111", b"00000000000000000000000000000000"),
	(b"11001101111100000011110111001011", b"01001110101111010110001000000100"), -- 2.09248e+09+-5.03823e+08=1.58866e+09
	(b"01001101000100100111000010000100", b"00000000000000000000000000000000"),
	(b"11001110100001000100101101110000", b"11001110011000111111101010111111"), -- 1.53553e+08+-1.10977e+09=-9.56215e+08
	(b"01001100110011000000000100100100", b"00000000000000000000000000000000"),
	(b"11001011111010010100000110101110", b"01001100100100011011000010111000"), -- 1.06957e+08+-3.05734e+07=7.63837e+07
	(b"11001110111000101100010110110100", b"00000000000000000000000000000000"),
	(b"11001110100111101110110011010011", b"11001111010000001101100101000100"), -- -1.9023e+09+-1.33316e+09=-3.23546e+09
	(b"11001101111011000010100110111001", b"00000000000000000000000000000000"),
	(b"11001101111010000010011110110100", b"11001110011010100010100010110110"), -- -4.9527e+08+-4.86865e+08=-9.82134e+08
	(b"11001110001100010100111010000000", b"00000000000000000000000000000000"),
	(b"11001110110011011111001100010111", b"11001111000100110100110100101100"), -- -7.43678e+08+-1.72763e+09=-2.47131e+09
	(b"11001110101101000001111110111100", b"00000000000000000000000000000000"),
	(b"11001110110111100000111000111001", b"11001111010010010001011011111010"), -- -1.51099e+09+-1.86274e+09=-3.37373e+09
	(b"11001101010011011111001000000000", b"00000000000000000000000000000000"),
	(b"01001101111100001001001000111111", b"01001101100010011001100100111111"), -- -2.15949e+08+5.04515e+08=2.88565e+08
	(b"01001110110000111001011010010000", b"00000000000000000000000000000000"),
	(b"01001110100111100010001000011110", b"01001111001100001101110001010111"), -- 1.64071e+09+1.32652e+09=2.96723e+09
	(b"01001101100000101100110111000111", b"00000000000000000000000000000000"),
	(b"01001110000100101100001011011000", b"01001110010101000010100110111100"), -- 2.74315e+08+6.15561e+08=8.89876e+08
	(b"11001110111100001010000101000111", b"00000000000000000000000000000000"),
	(b"01001110111010110110001100111110", b"11001100001001111100000100100000"), -- -2.01855e+09+1.97457e+09=-4.39758e+07
	(b"01001110101000010100101011010101", b"00000000000000000000000000000000"),
	(b"01001110111000011011011011001100", b"01001111010000011000000011010000"), -- 1.35302e+09+1.89343e+09=3.24644e+09
	(b"01001110100000010011011110110111", b"00000000000000000000000000000000"),
	(b"11001110111000100001101011100110", b"11001110010000011100011001011110"), -- 1.08396e+09+-1.89671e+09=-8.12751e+08
	(b"11001110110100101010111100011010", b"00000000000000000000000000000000"),
	(b"01001110101001101001001101000001", b"11001101101100000110111101100100"), -- -1.76735e+09+1.39733e+09=-3.70011e+08
	(b"11001110010000101110101011111101", b"00000000000000000000000000000000"),
	(b"11001110001101111111000001010101", b"11001110101111010110110110101001"), -- -8.17545e+08+-7.71495e+08=-1.58904e+09
	(b"01001101110001000100111110001101", b"00000000000000000000000000000000"),
	(b"01001110011010000110100111110011", b"01001110101001010100100011011101"), -- 4.11693e+08+9.74814e+08=1.38651e+09
	(b"11001101000100101011100011000000", b"00000000000000000000000000000000"),
	(b"01001101101010111011010111001111", b"01001101010001001011001011011110"), -- -1.53849e+08+3.60102e+08=2.06254e+08
	(b"11001110011010001001110111000000", b"00000000000000000000000000000000"),
	(b"11001110101110000010010000101100", b"11001111000101100011100110000110"), -- -9.75663e+08+-1.54469e+09=-2.52035e+09
	(b"11001110101000111000011101101010", b"00000000000000000000000000000000"),
	(b"11001110100011101101111010001110", b"11001111000110010011001011111100"), -- -1.37178e+09+-1.19848e+09=-2.57026e+09
	(b"11001110011000010010101010110101", b"00000000000000000000000000000000"),
	(b"01001110100110000011010111111010", b"01001101100111101000001001111110"), -- -9.44418e+08+1.27684e+09=3.32419e+08


	(x"3dcccccd", x"00000000"),
	(x"3dcccccd", x"3e4ccccd"),
	(x"c09ccccd", x"00000000"),
	(x"40a9999a", x"3ecccccd"),
	(x"40a9999a", x"00000000"),
	(x"c09ccccd", x"3ecccccd"),
	(x"c09ccccd", x"00000000"),
	(x"40a33333", x"3e4ccccd"),
	(x"40a33333", x"00000000"),
	(x"c09ccccd", x"3e4ccccd"),
	(x"c09ccccd", x"00000000"),
	(x"40a66666", x"3e99999a"),
	(x"40a66666", x"00000000"),
	(x"c09ccccd", x"3e99999a"),
	(x"c099999a", x"00000000"),
	(x"40a66666", x"3ecccccd"),
	(x"40a66666", x"00000000"),
	(x"c099999a", x"3ecccccd"),
	(x"653821cd", x"00000000"),
	(x"40a00033", x"653821cd"),
	(x"40200000", x"00000000"),
	(x"40a9999a", x"40f9999a"),
	(x"7f800000", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"7f800000", x"00000000"),
	(x"ff800000", x"7fffffff"),
	(x"ff800000", x"00000000"),
	(x"7f800000", x"7fffffff"),
	(x"ff800000", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"7f800000", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"7f800000", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"ff800000", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"ff800000", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"7fffffff", x"00000000"),
	(x"7f800000", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"7f800000", x"ffffffff"),
	(x"7fffffff", x"00000000"),
	(x"ff800000", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"ff800000", x"ffffffff"),
	(x"7fffffff", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"7fffffff", x"00000000"),
	(x"ffffffff", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"00000000", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"00000000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"00000000", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"80000000", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"80000000", x"ff800000"),
	(x"80000000", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"80000000", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"00000000", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"00000000", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"00000000", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"80000000", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"80000000", x"ffffffff"),
	(x"80000000", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"80000000", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"3f800000", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"3f800000", x"ff800000"),
	(x"3f800000", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"3f800000", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"bf800000", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"bf800000", x"ff800000"),
	(x"bf800000", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"bf800000", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"3f800000", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"3f800000", x"ffffffff"),
	(x"3f800000", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"3f800000", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"bf800000", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"bf800000", x"ffffffff"),
	(x"bf800000", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"bf800000", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"7bffffff", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"7bffffff", x"ff800000"),
	(x"7bffffff", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"7bffffff", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"fbffffff", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"fbffffff", x"ff800000"),
	(x"fbffffff", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"fbffffff", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"7bffffff", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"7bffffff", x"ffffffff"),
	(x"7bffffff", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"7bffffff", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"fbffffff", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"fbffffff", x"ffffffff"),
	(x"fbffffff", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"fbffffff", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"007fffff", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"007fffff", x"ff800000"),
	(x"007fffff", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"007fffff", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f800000", x"00000000"),
	(x"807fffff", x"7f800000"),
	(x"ff800000", x"00000000"),
	(x"807fffff", x"ff800000"),
	(x"807fffff", x"00000000"),
	(x"7f800000", x"7f800000"),
	(x"807fffff", x"00000000"),
	(x"ff800000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"007fffff", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"007fffff", x"ffffffff"),
	(x"007fffff", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"007fffff", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7fffffff", x"00000000"),
	(x"807fffff", x"7fffffff"),
	(x"ffffffff", x"00000000"),
	(x"807fffff", x"ffffffff"),
	(x"807fffff", x"00000000"),
	(x"7fffffff", x"7fffffff"),
	(x"807fffff", x"00000000"),
	(x"ffffffff", x"ffffffff"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"80000000", x"00000000"),
	(x"80000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"80000000", x"00000000"),
	(x"80000000", x"80000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7f000000", x"00000000"),
	(x"7f000000", x"7f800000"),
	(x"7f000000", x"00000000"),
	(x"ff000000", x"00000000"),
	(x"ff000000", x"00000000"),
	(x"7f000000", x"00000000"),
	(x"ff000000", x"00000000"),
	(x"ff000000", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"7e800000", x"00000000"),
	(x"7f000000", x"7f400000"),
	(x"7e800000", x"00000000"),
	(x"fe800000", x"00000000"),
	(x"fe800000", x"00000000"),
	(x"7e800000", x"00000000"),
	(x"ff000000", x"00000000"),
	(x"fe800000", x"ff400000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000001", x"00000000"),
	(x"00000001", x"00000002"),
	(x"00400000", x"00000000"),
	(x"00400000", x"00800000"),
	(x"7bffffff", x"00000000"),
	(x"7bffffff", x"7c7fffff"),
	(x"fbffffff", x"00000000"),
	(x"7bffffff", x"00000000"),
	(x"7bffffff", x"00000000"),
	(x"fbffffff", x"00000000"),
	(x"fbffffff", x"00000000"),
	(x"fbffffff", x"fc7fffff"),
	(x"7f7fffff", x"00000000"),
	(x"7f7fffff", x"7f800000"),
	(x"7f7fffff", x"00000000"),
	(x"ff7fffff", x"00000000"),
	(x"ff7fffff", x"00000000"),
	(x"7f7fffff", x"00000000"),
	(x"ff7fffff", x"00000000"),
	(x"ff7fffff", x"ff800000"),
	(x"bfe00000", x"00000000"),
	(x"40000000", x"3e800000"),
	(x"3fe00003", x"00000000"),
	(x"c0000007", x"be80002c"),
	(x"3fe00003", x"00000000"),
	(x"c0000005", x"be80001b"),
	(x"c0000005", x"00000000"),
	(x"3fe00003", x"be80001b"),
	(x"86844a7f", x"00000000"),
	(x"66844a7f", x"66844a7f"),
	(x"4004802b", x"00000000"),
	(x"3f04803d", x"4025a03a"),
	(x"55a5a03a", x"00000000"),
	(x"550da032", x"55ec7053"),
	(x"7f7fffff", x"00000000"),
	(x"7f7fffff", x"7f800000"),
	(x"80000001", x"00000000"),
	(x"80000001", x"80000002"),
	(x"ff7fffff", x"00000000"),
	(x"ff7fffff", x"ff800000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000"),
	(x"00000000", x"00000000")
	);



	---- Inf
	--		(x"7f800000", x"7f800000", x"7f800000"), -- inf + inf = inf
	--		(x"7f800000", x"ff800000", x"7fffffff"), -- inf + -inf = NaN	
	--		(x"ff800000", x"7f800000", x"7fffffff"), -- -inf + inf = NaN
	--		(x"ff800000", x"ff800000", x"ff800000"), -- -inf + -inf = -inf
	---- inf + NaN		
	--		(x"7f800000", x"7fffffff", x"7fffffff"), -- inf + NaN = NaN
	--		(x"7f800000", x"ffffffff", x"ffffffff"), -- inf + -NaN = -NaN
	--		(x"ff800000", x"7fffffff", x"7fffffff"), -- -inf + NaN = NaN
	--		(x"ff800000", x"ffffffff", x"ffffffff"), -- -inf + -NaN = -NaN
	---- NaN + inf
	--		(x"7fffffff", x"7f800000", x"7fffffff"), -- NaN + inf = NaN
	--		(x"ffffffff", x"7f800000", x"ffffffff"), -- -NaN + inf = -NaN
	--		(x"7fffffff", x"ff800000", x"7fffffff"), -- NaN + -inf = NaN
	--		(x"ffffffff", x"ff800000", x"ffffffff"), -- -NaN + -inf = -NaN		
	--
	---- TODO: Descobrir o que fazer com os NaN
	---- NaN
	--		(x"7fffffff", x"7fffffff", x"7fffffff"), -- NaN + NaN = NaN
	--		(x"7fffffff", x"ffffffff", x"7fffffff"), -- NaN + -NaN = NaN
	--		(x"ffffffff", x"7fffffff", x"7fffffff"), -- -NaN + NaN = NaN
	--		(x"ffffffff", x"ffffffff", x"ffffffff"), -- -NaN + -NaN = -NaN		
	---- Inf + 0
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7f800000", x"00000000", x"7f800000"), -- inf + 0 = inf
	--		(x"ff800000", x"00000000", x"ff800000"), -- -inf + 0 = -inf	
	--		(x"00000000", x"7f800000", x"7f800000"), -- 0 + inf = inf
	--		(x"00000000", x"ff800000", x"ff800000"), -- 0 + -inf = -inf
	---- inf + -0	
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7f800000", x"80000000", x"7f800000"), -- inf + -0 = inf
	--		(x"ff800000", x"80000000", x"ff800000"), -- -inf + -0 = -inf	
	--		(x"80000000", x"7f800000", x"7f800000"), -- -0 + inf = inf
	--		(x"80000000", x"ff800000", x"ff800000"), -- -0 + -inf = -inf
	---- NaN + 0
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"00000000", x"7fffffff"), -- NaN + 0 = NaN
	--		(x"ffffffff", x"00000000", x"ffffffff"), -- -NaN + 0 = -NaN	
	--		(x"00000000", x"7fffffff", x"7fffffff"), -- 0 + NaN = NaN
	--		(x"00000000", x"ffffffff", x"ffffffff"), -- 0 + -NaN = -NaN
	---- NaN + -0	
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"80000000", x"7fffffff"), -- NaN + -0 = NaN
	--		(x"ffffffff", x"80000000", x"ffffffff"), -- -NaN + -0 = -NaN	
	--		(x"80000000", x"7fffffff", x"7fffffff"), -- -0 + NaN = NaN
	--		(x"80000000", x"ffffffff", x"ffffffff"), -- -0 + -NaN = -NaN
	---- inf + 1		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7f800000", x"3f800000", x"7f800000"), -- inf + 1 = inf
	--		(x"ff800000", x"3f800000", x"ff800000"), -- -inf + 1 = -inf	
	--		(x"3f800000", x"7f800000", x"7f800000"), -- 1 + inf = inf
	--		(x"3f800000", x"ff800000", x"ff800000"), -- 1 + -inf = -inf
	---- inf + -1		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7f800000", x"bf800000", x"7f800000"), -- inf + -1 = inf
	--		(x"ff800000", x"bf800000", x"ff800000"), -- -inf + -1 = -inf	
	--		(x"bf800000", x"7f800000", x"7f800000"), -- -1 + inf = inf
	--		(x"bf800000", x"ff800000", x"ff800000"), -- -1 + -inf = -inf
	---- NaN + 1
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"3f800000", x"7fffffff"), -- NaN + 1 = NaN
	--		(x"ffffffff", x"3f800000", x"ffffffff"), -- -NaN + 1 = -NaN	
	--		(x"3f800000", x"7fffffff", x"7fffffff"), -- 1 + NaN = NaN
	--		(x"3f800000", x"ffffffff", x"ffffffff"), -- 1 + -NaN = -NaN
	---- Nan + -1		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"bf800000", x"7fffffff"), -- NaN + -1 = NaN
	--		(x"ffffffff", x"bf800000", x"ffffffff"), -- -NaN + -1 = -NaN	
	--		(x"bf800000", x"7fffffff", x"7fffffff"), -- -1 + NaN = NaN
	--		(x"bf800000", x"ffffffff", x"ffffffff"), -- -1 + -NaN = -NaN
	--		(x"00000000", x"00000000", x"00000000"),
	---- inf + 7bffffff		
	--		(x"7f800000", x"7bffffff", x"7f800000"), -- inf + 7bffffff = inf
	--		(x"ff800000", x"7bffffff", x"ff800000"), -- -inf + 7bffffff = -inf	
	--		(x"7bffffff", x"7f800000", x"7f800000"), -- 7bffffff + inf = inf
	--		(x"7bffffff", x"ff800000", x"ff800000"), -- 7bffffff + -inf = -inf
	---- inf + fbffffff		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7f800000", x"fbffffff", x"7f800000"), -- inf + -fbffffff = inf
	--		(x"ff800000", x"fbffffff", x"ff800000"), -- -inf + -fbffffff = -inf	
	--		(x"fbffffff", x"7f800000", x"7f800000"), -- -fbffffff + inf = inf
	--		(x"fbffffff", x"ff800000", x"ff800000"), -- -fbffffff + -inf = -inf
	---- NaN + 7bffffff
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"7bffffff", x"7fffffff"), -- NaN + 7bffffff = NaN
	--		(x"ffffffff", x"7bffffff", x"ffffffff"), -- -NaN + 7bffffff = -NaN	
	--		(x"7bffffff", x"7fffffff", x"7fffffff"), -- 7bffffff + NaN = NaN
	--		(x"7bffffff", x"ffffffff", x"ffffffff"), -- 7bffffff + -NaN = -NaN
	---- Nan + fbffffff		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"fbffffff", x"7fffffff"), -- NaN + fbffffff = NaN
	--		(x"ffffffff", x"fbffffff", x"ffffffff"), -- -NaN + fbffffff = -NaN	
	--		(x"fbffffff", x"7fffffff", x"7fffffff"), -- fbffffff + NaN = NaN
	--		(x"fbffffff", x"ffffffff", x"ffffffff"), -- fbffffff + -NaN = -NaN
	--		(x"00000000", x"00000000", x"00000000"),
	---- inf + 007fffff		
	--		(x"7f800000", x"007fffff", x"7f800000"), -- inf + 007fffff = inf
	--		(x"ff800000", x"007fffff", x"ff800000"), -- -inf + 007fffff = -inf	
	--		(x"007fffff", x"7f800000", x"7f800000"), -- 007fffff + inf = inf
	--		(x"007fffff", x"ff800000", x"ff800000"), -- 007fffff + -inf = -inf
	---- inf + 807fffff		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7f800000", x"807fffff", x"7f800000"), -- inf + 807fffff = inf
	--		(x"ff800000", x"807fffff", x"ff800000"), -- -inf + 807fffff = -inf	
	--		(x"807fffff", x"7f800000", x"7f800000"), -- 807fffff + inf = inf
	--		(x"807fffff", x"ff800000", x"ff800000"), -- 807fffff + -inf = -inf
	---- NaN + 007fffff
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"007fffff", x"7fffffff"), -- NaN + 007fffff = NaN
	--		(x"ffffffff", x"007fffff", x"ffffffff"), -- -NaN + 007fffff = -NaN	
	--		(x"007fffff", x"7fffffff", x"7fffffff"), -- 007fffff + NaN = NaN
	--		(x"007fffff", x"ffffffff", x"ffffffff"), -- 007fffff + -NaN = -NaN
	---- Nan + 807fffff		
	--		(x"00000000", x"00000000", x"00000000"),
	--		(x"7fffffff", x"807fffff", x"7fffffff"), -- NaN + 807fffff = NaN
	--		(x"ffffffff", x"807fffff", x"ffffffff"), -- -NaN + 807fffff = -NaN	
	--		(x"807fffff", x"7fffffff", x"7fffffff"), -- 807fffff + NaN = NaN
	--		(x"807fffff", x"ffffffff", x"ffffffff"), -- 807fffff + -NaN = -NaN
	--		(x"00000000", x"00000000", x"00000000"),
	---- 0 + -0		
	--		(x"00000000", x"00000000", x"00000000"), -- 0 + 0 = 0
	--		(x"00000000", x"80000000", x"00000000"), -- 0 + -0 = 0
	--		(x"80000000", x"00000000", x"00000000"), -- -0 + 0 = 0
	--		(x"80000000", x"80000000", x"80000000"), -- -0 + -0 = -0
	--		(x"00000000", x"00000000", x"00000000"),
	--
	---- Overflow
	--		(x"7f000000", x"7f000000", x"7f800000"), -- 7f000000 + 7f000000 = inf
	--		(x"7f000000", x"ff000000", x"00000000"), -- 7f000000 + ff000000 = 0
	--		(x"ff000000", x"7f000000", x"00000000"), -- ff000000 + 7f000000 = 0
	--		(x"ff000000", x"ff000000", x"ff800000"), -- ff000000 + ff000000 = -inf
	--		(x"00000000", x"00000000", x"00000000"),
	--		
	--		(x"7e800000", x"7f000000", x"7f400000"), -- 7e800000 + 7f000000 = 7f400000 # não é overflow
	--		(x"7e800000", x"fe800000", x"00000000"), -- 7e800000 + fe800000 = 0
	--		(x"fe800000", x"7e800000", x"00000000"), -- fe800000 + 7e800000 = 0
	--		(x"ff000000", x"fe800000", x"ff400000"), -- ff000000 + fe800000 = -inf	   # não é overflow
	--		(x"00000000", x"00000000", x"00000000"),
	--
	---- Denormalized
	--		(x"00000001", x"00000001", x"00000002"), -- 00000001 + 00000001 = 00000002
	--		(x"00400000", x"00400000", x"00800000"), -- 00400000 + 00400000 = 00800000 
	---- Round
	--		(x"7bffffff", x"7bffffff", x"7c7fffff"), -- 7bffffff + 7bffffff = 7c7fffff
	--		(x"fbffffff", x"7bffffff", x"00000000"), -- fbffffff + 7bffffff = 0
	--		(x"7bffffff", x"fbffffff", x"00000000"), -- 7bffffff + fbffffff = 0
	--		(x"fbffffff", x"fbffffff", x"ff800000"), -- fbffffff + fbffffff = -inf
	--		
	--		(x"7f7fffff", x"7f7fffff", x"7f800000"), -- 7f7fffff + 7f7fffff = inf
	--		(x"7f7fffff", x"ff7fffff", x"00000000"), -- 7f7fffff + ff7fffff = 0
	--		(x"ff7fffff", x"7f7fffff", x"00000000"), -- ff7fffff + 7f7fffff = 0
	--		(x"ff7fffff", x"ff7fffff", x"ff800000"), -- ff7fffff + ff7fffff = -inf
	--		
	--		(x"bfe00000", x"40000000", x"3e800000"),
	--		(x"3fe00003", x"c0000007", x"be80002c"),
	--		(x"3fe00003", x"c0000005", x"be80001b"),
	--		(x"86844a7f", x"66844a7f", x"66844a7f"), -- 4.9762344E-35 	3.123633E23
	--		(x"4004802b", x"3f04803d", x"4025a03a"), -- 2.0703228 		0.51758176 --		2.5879045
	--		(x"55a5a03a", x"550da032", x"55ec7053"), -- 9.7324483E12 	2.27634483E13 	3.24958966E13
	--		(x"7f7fffff", x"7f7fffff", x"00000000"),
	--		(x"80000001", x"80000001", x"00000000"),
	--		(x"ff7fffff", x"ff7fffff", x"00000000"),
	--		(x"00000000", x"00000000", x"00000000")

	begin
	--	clock <= not clock after 200 NS;

	reset <= '1', '0' after 250 NS;

	clk: process
	begin
		clock <= '0';
		wait for 200 ns;
		clock <= '1';
		wait for 200 ns;
	end process clk;	

	sel: process
	begin
		wait until rising_edge(clock);
		sela <= '1';
		selb <= '0';
		wait until rising_edge(clock);
		sela <= '0';
		selb <= '1';
	end process;

	--	rst: process
	--	begin
	--		reset <= '0';
	--		wait for 250 ns;
	--		reset <= '1';
	--	end process rst;	

	--	f2 <= "00111111111000000000000000000000" after 500 NS;
	--	f1 <= "11000000000000000000000000000000" after 500 NS;

	Gera_entradas: process
	variable v : entrada;
	begin

		for i in test_vector'range loop
			wait until rising_edge(clock);
			v := test_vector(i);
			AB_in <= v.a;
			f3_tmp <= v.b;
			f3_tmp2 <= f3_tmp;
			f3 <= f3_tmp2;
		end loop;

		--	f2 <= "10111111111000000000000000000000";
		--	f1 <= "01000000000000000000000000000000";
		--	f2 <= "00111111111000000000000000000011" after 950 NS;
		--	f1 <= "11000000000000000000000000000111" after 950 NS;
		--	f2 <= "00111111111000000000000000000011" after 1150 NS;
		--	f1 <= "11000000000000000000000000000101" after 1150 NS;
	end process Gera_entradas;


	process (res, f3, selb)
	begin
		if ((res = f3) or (selb = '0')) then
			ok <= '1';
		else
			ok <= '0';
		end if;
		if (res(30 downto 23) = f3(30 downto 23) or (selb='0')) then
			ok_exp <= '1';
		else
			ok_exp <= '0';
		end if;
	end process;

		--	segura1: process
		--	begin
		--		wait until rising_edge(clock);
		--		auxv1 <= f3;
		--	end process segura1;
		--	
		--	segura2: process
		--	begin
		--		wait until rising_edge(clock);
		--		auxv2 <= auxv1;
		--	end process segura2;
		--	
	--	compara_resultados: process(auxv2, res)
		--	begin
		--		if (auxv2 = res) then
		--			aux <= '1';
		--		else
		--			aux <= '0';
		--		end if;
		--	end process compara_resultados;
		--	ok <= aux;

		--selb <= not sela;

	A: entity work.somador port map (AB_in, clock, reset, wt_in, sela, selb, selc, res, pronto, wt_out);
end arch_somador;
